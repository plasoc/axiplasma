library ieee;
use ieee.std_logic_1164.all;

package ram_pack is

	constant cpu_width : integer := 32;
	constant ram_size : integer := 16384;
	subtype word_type is std_logic_vector(cpu_width-1 downto 0);
	type ram_type is array(0 to ram_size-1) of word_type;
	function load_hex return ram_type;

end package;

package body ram_pack is

	function load_hex return ram_type is
		variable ram_buffer : ram_type := (others=>(others=>'0'));
	begin
		ram_buffer(0) := X"3C1C0101";
		ram_buffer(1) := X"279CD590";
		ram_buffer(2) := X"3C050100";
		ram_buffer(3) := X"24A55598";
		ram_buffer(4) := X"3C040101";
		ram_buffer(5) := X"248459BC";
		ram_buffer(6) := X"3C1D0101";
		ram_buffer(7) := X"27BD58E8";
		ram_buffer(8) := X"ACA00000";
		ram_buffer(9) := X"00A4182A";
		ram_buffer(10) := X"1460FFFD";
		ram_buffer(11) := X"24A50004";
		ram_buffer(12) := X"0C40007C";
		ram_buffer(13) := X"00000000";
		ram_buffer(14) := X"0840000E";
		ram_buffer(15) := X"23BDFF98";
		ram_buffer(16) := X"AFA10010";
		ram_buffer(17) := X"AFA20014";
		ram_buffer(18) := X"AFA30018";
		ram_buffer(19) := X"AFA4001C";
		ram_buffer(20) := X"AFA50020";
		ram_buffer(21) := X"AFA60024";
		ram_buffer(22) := X"AFA70028";
		ram_buffer(23) := X"AFA8002C";
		ram_buffer(24) := X"AFA90030";
		ram_buffer(25) := X"AFAA0034";
		ram_buffer(26) := X"AFAB0038";
		ram_buffer(27) := X"AFAC003C";
		ram_buffer(28) := X"AFAD0040";
		ram_buffer(29) := X"AFAE0044";
		ram_buffer(30) := X"AFAF0048";
		ram_buffer(31) := X"AFB8004C";
		ram_buffer(32) := X"AFB90050";
		ram_buffer(33) := X"AFBF0054";
		ram_buffer(34) := X"401A7000";
		ram_buffer(35) := X"235AFFFC";
		ram_buffer(36) := X"AFBA0058";
		ram_buffer(37) := X"0000D810";
		ram_buffer(38) := X"AFBB005C";
		ram_buffer(39) := X"0000D812";
		ram_buffer(40) := X"AFBB0060";
		ram_buffer(41) := X"0C4012B2";
		ram_buffer(42) := X"23A50000";
		ram_buffer(43) := X"8FA10010";
		ram_buffer(44) := X"8FA20014";
		ram_buffer(45) := X"8FA30018";
		ram_buffer(46) := X"8FA4001C";
		ram_buffer(47) := X"8FA50020";
		ram_buffer(48) := X"8FA60024";
		ram_buffer(49) := X"8FA70028";
		ram_buffer(50) := X"8FA8002C";
		ram_buffer(51) := X"8FA90030";
		ram_buffer(52) := X"8FAA0034";
		ram_buffer(53) := X"8FAB0038";
		ram_buffer(54) := X"8FAC003C";
		ram_buffer(55) := X"8FAD0040";
		ram_buffer(56) := X"8FAE0044";
		ram_buffer(57) := X"8FAF0048";
		ram_buffer(58) := X"8FB8004C";
		ram_buffer(59) := X"8FB90050";
		ram_buffer(60) := X"8FBF0054";
		ram_buffer(61) := X"8FBA0058";
		ram_buffer(62) := X"8FBB005C";
		ram_buffer(63) := X"03600011";
		ram_buffer(64) := X"8FBB0060";
		ram_buffer(65) := X"03600013";
		ram_buffer(66) := X"23BD0068";
		ram_buffer(67) := X"341B0001";
		ram_buffer(68) := X"03400008";
		ram_buffer(69) := X"409B6000";
		ram_buffer(70) := X"40026000";
		ram_buffer(71) := X"03E00008";
		ram_buffer(72) := X"40846000";
		ram_buffer(73) := X"3C050100";
		ram_buffer(74) := X"24A50150";
		ram_buffer(75) := X"8CA60000";
		ram_buffer(76) := X"AC06003C";
		ram_buffer(77) := X"8CA60004";
		ram_buffer(78) := X"AC060040";
		ram_buffer(79) := X"8CA60008";
		ram_buffer(80) := X"AC060044";
		ram_buffer(81) := X"8CA6000C";
		ram_buffer(82) := X"03E00008";
		ram_buffer(83) := X"AC060048";
		ram_buffer(84) := X"3C1A0100";
		ram_buffer(85) := X"375A003C";
		ram_buffer(86) := X"03400008";
		ram_buffer(87) := X"00000000";
		ram_buffer(88) := X"AC900000";
		ram_buffer(89) := X"AC910004";
		ram_buffer(90) := X"AC920008";
		ram_buffer(91) := X"AC93000C";
		ram_buffer(92) := X"AC940010";
		ram_buffer(93) := X"AC950014";
		ram_buffer(94) := X"AC960018";
		ram_buffer(95) := X"AC97001C";
		ram_buffer(96) := X"AC9E0020";
		ram_buffer(97) := X"AC9C0024";
		ram_buffer(98) := X"AC9D0028";
		ram_buffer(99) := X"AC9F002C";
		ram_buffer(100) := X"03E00008";
		ram_buffer(101) := X"34020000";
		ram_buffer(102) := X"8C900000";
		ram_buffer(103) := X"8C910004";
		ram_buffer(104) := X"8C920008";
		ram_buffer(105) := X"8C93000C";
		ram_buffer(106) := X"8C940010";
		ram_buffer(107) := X"8C950014";
		ram_buffer(108) := X"8C960018";
		ram_buffer(109) := X"8C97001C";
		ram_buffer(110) := X"8C9E0020";
		ram_buffer(111) := X"8C9C0024";
		ram_buffer(112) := X"8C9D0028";
		ram_buffer(113) := X"8C9F002C";
		ram_buffer(114) := X"03E00008";
		ram_buffer(115) := X"34A20000";
		ram_buffer(116) := X"00850019";
		ram_buffer(117) := X"00001012";
		ram_buffer(118) := X"00002010";
		ram_buffer(119) := X"03E00008";
		ram_buffer(120) := X"ACC40000";
		ram_buffer(121) := X"0000000C";
		ram_buffer(122) := X"03E00008";
		ram_buffer(123) := X"00000000";
		ram_buffer(124) := X"3C040100";
		ram_buffer(125) := X"27BDFFE8";
		ram_buffer(126) := X"AFBF0014";
		ram_buffer(127) := X"0C40028D";
		ram_buffer(128) := X"248404AC";
		ram_buffer(129) := X"8FBF0014";
		ram_buffer(130) := X"00001025";
		ram_buffer(131) := X"03E00008";
		ram_buffer(132) := X"27BD0018";
		ram_buffer(133) := X"2082FF78";
		ram_buffer(134) := X"AC450078";
		ram_buffer(135) := X"03E00008";
		ram_buffer(136) := X"AC46001C";
		ram_buffer(137) := X"3C1A0100";
		ram_buffer(138) := X"375A5600";
		ram_buffer(139) := X"8F5B0000";
		ram_buffer(140) := X"AF400000";
		ram_buffer(141) := X"23BDFF78";
		ram_buffer(142) := X"AFA10010";
		ram_buffer(143) := X"AFA20014";
		ram_buffer(144) := X"AFA30018";
		ram_buffer(145) := X"AFA4001C";
		ram_buffer(146) := X"AFA50020";
		ram_buffer(147) := X"AFA60024";
		ram_buffer(148) := X"AFA70028";
		ram_buffer(149) := X"AFA8002C";
		ram_buffer(150) := X"AFA90030";
		ram_buffer(151) := X"AFAA0034";
		ram_buffer(152) := X"AFAB0038";
		ram_buffer(153) := X"AFAC003C";
		ram_buffer(154) := X"AFAD0040";
		ram_buffer(155) := X"AFAE0044";
		ram_buffer(156) := X"AFAF0048";
		ram_buffer(157) := X"AFB0004C";
		ram_buffer(158) := X"AFB10050";
		ram_buffer(159) := X"AFB20054";
		ram_buffer(160) := X"AFB30058";
		ram_buffer(161) := X"AFB4005C";
		ram_buffer(162) := X"AFB50060";
		ram_buffer(163) := X"AFB60064";
		ram_buffer(164) := X"AFB70068";
		ram_buffer(165) := X"AFB8006C";
		ram_buffer(166) := X"AFB90070";
		ram_buffer(167) := X"AFBF0074";
		ram_buffer(168) := X"401A7000";
		ram_buffer(169) := X"17600003";
		ram_buffer(170) := X"235AFFFC";
		ram_buffer(171) := X"084000AE";
		ram_buffer(172) := X"00000000";
		ram_buffer(173) := X"235A0004";
		ram_buffer(174) := X"AFBA0078";
		ram_buffer(175) := X"0000D810";
		ram_buffer(176) := X"AFBB007C";
		ram_buffer(177) := X"0000D812";
		ram_buffer(178) := X"AFBB0080";
		ram_buffer(179) := X"3C1A0100";
		ram_buffer(180) := X"375A55A8";
		ram_buffer(181) := X"8F5A0000";
		ram_buffer(182) := X"AF5D0000";
		ram_buffer(183) := X"3C1A0101";
		ram_buffer(184) := X"375A5700";
		ram_buffer(185) := X"8F5D0000";
		ram_buffer(186) := X"0C40023C";
		ram_buffer(187) := X"00000000";
		ram_buffer(188) := X"3C1A0101";
		ram_buffer(189) := X"375A5700";
		ram_buffer(190) := X"AF5D0000";
		ram_buffer(191) := X"3C1A0100";
		ram_buffer(192) := X"375A55A8";
		ram_buffer(193) := X"8F5A0000";
		ram_buffer(194) := X"8F5D0000";
		ram_buffer(195) := X"8FA10010";
		ram_buffer(196) := X"8FA20014";
		ram_buffer(197) := X"8FA30018";
		ram_buffer(198) := X"8FA4001C";
		ram_buffer(199) := X"8FA50020";
		ram_buffer(200) := X"8FA60024";
		ram_buffer(201) := X"8FA70028";
		ram_buffer(202) := X"8FA8002C";
		ram_buffer(203) := X"8FA90030";
		ram_buffer(204) := X"8FAA0034";
		ram_buffer(205) := X"8FAB0038";
		ram_buffer(206) := X"8FAC003C";
		ram_buffer(207) := X"8FAD0040";
		ram_buffer(208) := X"8FAE0044";
		ram_buffer(209) := X"8FAF0048";
		ram_buffer(210) := X"8FB0004C";
		ram_buffer(211) := X"8FB10050";
		ram_buffer(212) := X"8FB20054";
		ram_buffer(213) := X"8FB30058";
		ram_buffer(214) := X"8FB4005C";
		ram_buffer(215) := X"8FB50060";
		ram_buffer(216) := X"8FB60064";
		ram_buffer(217) := X"8FB70068";
		ram_buffer(218) := X"8FB8006C";
		ram_buffer(219) := X"8FB90070";
		ram_buffer(220) := X"8FBF0074";
		ram_buffer(221) := X"8FBA0078";
		ram_buffer(222) := X"8FBB007C";
		ram_buffer(223) := X"03600011";
		ram_buffer(224) := X"8FBB0080";
		ram_buffer(225) := X"03600013";
		ram_buffer(226) := X"23BD0088";
		ram_buffer(227) := X"341B0001";
		ram_buffer(228) := X"03400008";
		ram_buffer(229) := X"409B6000";
		ram_buffer(230) := X"00000000";
		ram_buffer(231) := X"3C080100";
		ram_buffer(232) := X"250803C8";
		ram_buffer(233) := X"8D090000";
		ram_buffer(234) := X"AC09003C";
		ram_buffer(235) := X"8D090004";
		ram_buffer(236) := X"AC090040";
		ram_buffer(237) := X"8D090008";
		ram_buffer(238) := X"AC090044";
		ram_buffer(239) := X"8D09000C";
		ram_buffer(240) := X"03E00008";
		ram_buffer(241) := X"AC090048";
		ram_buffer(242) := X"3C1A0100";
		ram_buffer(243) := X"375A0224";
		ram_buffer(244) := X"03400008";
		ram_buffer(245) := X"00000000";
		ram_buffer(246) := X"3C1A0101";
		ram_buffer(247) := X"375A5700";
		ram_buffer(248) := X"AF5D0000";
		ram_buffer(249) := X"3C1A0100";
		ram_buffer(250) := X"375A55A8";
		ram_buffer(251) := X"8F5A0000";
		ram_buffer(252) := X"8F5D0000";
		ram_buffer(253) := X"8FA10010";
		ram_buffer(254) := X"8FA20014";
		ram_buffer(255) := X"8FA30018";
		ram_buffer(256) := X"8FA4001C";
		ram_buffer(257) := X"8FA50020";
		ram_buffer(258) := X"8FA60024";
		ram_buffer(259) := X"8FA70028";
		ram_buffer(260) := X"8FA8002C";
		ram_buffer(261) := X"8FA90030";
		ram_buffer(262) := X"8FAA0034";
		ram_buffer(263) := X"8FAB0038";
		ram_buffer(264) := X"8FAC003C";
		ram_buffer(265) := X"8FAD0040";
		ram_buffer(266) := X"8FAE0044";
		ram_buffer(267) := X"8FAF0048";
		ram_buffer(268) := X"8FB0004C";
		ram_buffer(269) := X"8FB10050";
		ram_buffer(270) := X"8FB20054";
		ram_buffer(271) := X"8FB30058";
		ram_buffer(272) := X"8FB4005C";
		ram_buffer(273) := X"8FB50060";
		ram_buffer(274) := X"8FB60064";
		ram_buffer(275) := X"8FB70068";
		ram_buffer(276) := X"8FB8006C";
		ram_buffer(277) := X"8FB90070";
		ram_buffer(278) := X"8FBF0074";
		ram_buffer(279) := X"8FBA0078";
		ram_buffer(280) := X"8FBB007C";
		ram_buffer(281) := X"03600011";
		ram_buffer(282) := X"8FBB0080";
		ram_buffer(283) := X"03600013";
		ram_buffer(284) := X"23BD0088";
		ram_buffer(285) := X"341B0001";
		ram_buffer(286) := X"03400008";
		ram_buffer(287) := X"409B6000";
		ram_buffer(288) := X"40806000";
		ram_buffer(289) := X"20090001";
		ram_buffer(290) := X"3C080100";
		ram_buffer(291) := X"35085600";
		ram_buffer(292) := X"AD090000";
		ram_buffer(293) := X"3C080100";
		ram_buffer(294) := X"350855E4";
		ram_buffer(295) := X"AD090000";
		ram_buffer(296) := X"0000000C";
		ram_buffer(297) := X"03E00008";
		ram_buffer(298) := X"00000000";
		ram_buffer(299) := X"3C060100";
		ram_buffer(300) := X"27BDFFE8";
		ram_buffer(301) := X"24C60544";
		ram_buffer(302) := X"2405001E";
		ram_buffer(303) := X"AFBF0014";
		ram_buffer(304) := X"0C4002BF";
		ram_buffer(305) := X"00002025";
		ram_buffer(306) := X"3C060100";
		ram_buffer(307) := X"24C60580";
		ram_buffer(308) := X"24050018";
		ram_buffer(309) := X"0C4002BF";
		ram_buffer(310) := X"24040001";
		ram_buffer(311) := X"3C060100";
		ram_buffer(312) := X"24C605CC";
		ram_buffer(313) := X"24050012";
		ram_buffer(314) := X"0C4002BF";
		ram_buffer(315) := X"24040002";
		ram_buffer(316) := X"3C060100";
		ram_buffer(317) := X"24C60618";
		ram_buffer(318) := X"2405000C";
		ram_buffer(319) := X"0C4002BF";
		ram_buffer(320) := X"24040003";
		ram_buffer(321) := X"3C060100";
		ram_buffer(322) := X"24C60664";
		ram_buffer(323) := X"24050006";
		ram_buffer(324) := X"0C4002BF";
		ram_buffer(325) := X"24040004";
		ram_buffer(326) := X"0C4002DF";
		ram_buffer(327) := X"00002025";
		ram_buffer(328) := X"3C060100";
		ram_buffer(329) := X"24040005";
		ram_buffer(330) := X"24C606AC";
		ram_buffer(331) := X"0C4002BF";
		ram_buffer(332) := X"24050002";
		ram_buffer(333) := X"8FBF0014";
		ram_buffer(334) := X"24040005";
		ram_buffer(335) := X"084002DF";
		ram_buffer(336) := X"27BD0018";
		ram_buffer(337) := X"27BDFFE0";
		ram_buffer(338) := X"AFB10018";
		ram_buffer(339) := X"AFB00014";
		ram_buffer(340) := X"AFBF001C";
		ram_buffer(341) := X"3C1044A2";
		ram_buffer(342) := X"2411000F";
		ram_buffer(343) := X"0C4002DF";
		ram_buffer(344) := X"24040001";
		ram_buffer(345) := X"8F828084";
		ram_buffer(346) := X"00000000";
		ram_buffer(347) := X"24420001";
		ram_buffer(348) := X"AF828084";
		ram_buffer(349) := X"AE110008";
		ram_buffer(350) := X"1000FFF8";
		ram_buffer(351) := X"00000000";
		ram_buffer(352) := X"27BDFFE0";
		ram_buffer(353) := X"24040001";
		ram_buffer(354) := X"AFB10018";
		ram_buffer(355) := X"AFB00014";
		ram_buffer(356) := X"AFBF001C";
		ram_buffer(357) := X"0C4002F5";
		ram_buffer(358) := X"3C1044A2";
		ram_buffer(359) := X"2411001F";
		ram_buffer(360) := X"0C4002DF";
		ram_buffer(361) := X"24040002";
		ram_buffer(362) := X"8F828080";
		ram_buffer(363) := X"24040001";
		ram_buffer(364) := X"24420001";
		ram_buffer(365) := X"AF828080";
		ram_buffer(366) := X"AE110008";
		ram_buffer(367) := X"0C4002F5";
		ram_buffer(368) := X"00000000";
		ram_buffer(369) := X"1000FFF6";
		ram_buffer(370) := X"00000000";
		ram_buffer(371) := X"27BDFFE0";
		ram_buffer(372) := X"24040002";
		ram_buffer(373) := X"AFB10018";
		ram_buffer(374) := X"AFB00014";
		ram_buffer(375) := X"AFBF001C";
		ram_buffer(376) := X"0C4002F5";
		ram_buffer(377) := X"3C1044A2";
		ram_buffer(378) := X"2411002F";
		ram_buffer(379) := X"0C4002DF";
		ram_buffer(380) := X"24040003";
		ram_buffer(381) := X"8F82807C";
		ram_buffer(382) := X"24040002";
		ram_buffer(383) := X"24420001";
		ram_buffer(384) := X"AF82807C";
		ram_buffer(385) := X"AE110008";
		ram_buffer(386) := X"0C4002F5";
		ram_buffer(387) := X"00000000";
		ram_buffer(388) := X"1000FFF6";
		ram_buffer(389) := X"00000000";
		ram_buffer(390) := X"27BDFFE0";
		ram_buffer(391) := X"24040003";
		ram_buffer(392) := X"AFB10018";
		ram_buffer(393) := X"AFB00014";
		ram_buffer(394) := X"AFBF001C";
		ram_buffer(395) := X"0C4002F5";
		ram_buffer(396) := X"3C1044A2";
		ram_buffer(397) := X"2411003F";
		ram_buffer(398) := X"0C4002DF";
		ram_buffer(399) := X"24040004";
		ram_buffer(400) := X"8F828074";
		ram_buffer(401) := X"24040003";
		ram_buffer(402) := X"24420001";
		ram_buffer(403) := X"AF828074";
		ram_buffer(404) := X"AE110008";
		ram_buffer(405) := X"0C4002F5";
		ram_buffer(406) := X"00000000";
		ram_buffer(407) := X"1000FFF6";
		ram_buffer(408) := X"00000000";
		ram_buffer(409) := X"27BDFFE0";
		ram_buffer(410) := X"24040004";
		ram_buffer(411) := X"AFB00014";
		ram_buffer(412) := X"3C1044A2";
		ram_buffer(413) := X"AFB10018";
		ram_buffer(414) := X"AFBF001C";
		ram_buffer(415) := X"0C4002F5";
		ram_buffer(416) := X"26100008";
		ram_buffer(417) := X"2411004F";
		ram_buffer(418) := X"8F828078";
		ram_buffer(419) := X"24040004";
		ram_buffer(420) := X"24420001";
		ram_buffer(421) := X"AF828078";
		ram_buffer(422) := X"AE110000";
		ram_buffer(423) := X"0C4002F5";
		ram_buffer(424) := X"00000000";
		ram_buffer(425) := X"1000FFF8";
		ram_buffer(426) := X"00000000";
		ram_buffer(427) := X"27BDFFD0";
		ram_buffer(428) := X"AFB50024";
		ram_buffer(429) := X"AFB40020";
		ram_buffer(430) := X"AFB20018";
		ram_buffer(431) := X"AFB10014";
		ram_buffer(432) := X"3C140100";
		ram_buffer(433) := X"3C150100";
		ram_buffer(434) := X"3C120100";
		ram_buffer(435) := X"3C110100";
		ram_buffer(436) := X"AFB60028";
		ram_buffer(437) := X"AFB3001C";
		ram_buffer(438) := X"AFBF002C";
		ram_buffer(439) := X"AFB00010";
		ram_buffer(440) := X"0000B025";
		ram_buffer(441) := X"00009825";
		ram_buffer(442) := X"269452F4";
		ram_buffer(443) := X"26B5533C";
		ram_buffer(444) := X"265253AC";
		ram_buffer(445) := X"263153E0";
		ram_buffer(446) := X"2404001E";
		ram_buffer(447) := X"0C400304";
		ram_buffer(448) := X"2673001E";
		ram_buffer(449) := X"02602825";
		ram_buffer(450) := X"0C4004DC";
		ram_buffer(451) := X"02802025";
		ram_buffer(452) := X"8F908084";
		ram_buffer(453) := X"8F858080";
		ram_buffer(454) := X"8F84807C";
		ram_buffer(455) := X"02058021";
		ram_buffer(456) := X"8F838074";
		ram_buffer(457) := X"02048021";
		ram_buffer(458) := X"8F828078";
		ram_buffer(459) := X"02038021";
		ram_buffer(460) := X"02028021";
		ram_buffer(461) := X"24020005";
		ram_buffer(462) := X"14400002";
		ram_buffer(463) := X"0202001B";
		ram_buffer(464) := X"0007000D";
		ram_buffer(465) := X"8F848084";
		ram_buffer(466) := X"00001012";
		ram_buffer(467) := X"2443FFFF";
		ram_buffer(468) := X"0083202B";
		ram_buffer(469) := X"1480002E";
		ram_buffer(470) := X"00000000";
		ram_buffer(471) := X"8F848084";
		ram_buffer(472) := X"24420001";
		ram_buffer(473) := X"0044202B";
		ram_buffer(474) := X"14800029";
		ram_buffer(475) := X"00000000";
		ram_buffer(476) := X"8F848080";
		ram_buffer(477) := X"00000000";
		ram_buffer(478) := X"0083202B";
		ram_buffer(479) := X"14800024";
		ram_buffer(480) := X"00000000";
		ram_buffer(481) := X"8F848080";
		ram_buffer(482) := X"00000000";
		ram_buffer(483) := X"0044202B";
		ram_buffer(484) := X"1480001F";
		ram_buffer(485) := X"00000000";
		ram_buffer(486) := X"8F84807C";
		ram_buffer(487) := X"00000000";
		ram_buffer(488) := X"0083202B";
		ram_buffer(489) := X"1480001A";
		ram_buffer(490) := X"00000000";
		ram_buffer(491) := X"8F84807C";
		ram_buffer(492) := X"00000000";
		ram_buffer(493) := X"0044202B";
		ram_buffer(494) := X"14800015";
		ram_buffer(495) := X"00000000";
		ram_buffer(496) := X"8F848074";
		ram_buffer(497) := X"00000000";
		ram_buffer(498) := X"0083202B";
		ram_buffer(499) := X"14800010";
		ram_buffer(500) := X"00000000";
		ram_buffer(501) := X"8F848074";
		ram_buffer(502) := X"00000000";
		ram_buffer(503) := X"0044202B";
		ram_buffer(504) := X"1480000B";
		ram_buffer(505) := X"00000000";
		ram_buffer(506) := X"8F848078";
		ram_buffer(507) := X"00000000";
		ram_buffer(508) := X"0083182B";
		ram_buffer(509) := X"14600006";
		ram_buffer(510) := X"00000000";
		ram_buffer(511) := X"8F838078";
		ram_buffer(512) := X"00000000";
		ram_buffer(513) := X"0043102B";
		ram_buffer(514) := X"10400003";
		ram_buffer(515) := X"00000000";
		ram_buffer(516) := X"0C4004DC";
		ram_buffer(517) := X"02A02025";
		ram_buffer(518) := X"8F858084";
		ram_buffer(519) := X"0C4004DC";
		ram_buffer(520) := X"02402025";
		ram_buffer(521) := X"8F858080";
		ram_buffer(522) := X"0C4004DC";
		ram_buffer(523) := X"02202025";
		ram_buffer(524) := X"8F85807C";
		ram_buffer(525) := X"3C040100";
		ram_buffer(526) := X"0C4004DC";
		ram_buffer(527) := X"24845414";
		ram_buffer(528) := X"8F858074";
		ram_buffer(529) := X"3C040100";
		ram_buffer(530) := X"0C4004DC";
		ram_buffer(531) := X"24845448";
		ram_buffer(532) := X"8F858078";
		ram_buffer(533) := X"3C040100";
		ram_buffer(534) := X"0C4004DC";
		ram_buffer(535) := X"2484547C";
		ram_buffer(536) := X"3C040100";
		ram_buffer(537) := X"02162823";
		ram_buffer(538) := X"0C4004DC";
		ram_buffer(539) := X"248454B0";
		ram_buffer(540) := X"1000FFA1";
		ram_buffer(541) := X"0200B025";
		ram_buffer(542) := X"8F838094";
		ram_buffer(543) := X"00000000";
		ram_buffer(544) := X"8C620000";
		ram_buffer(545) := X"00000000";
		ram_buffer(546) := X"30420002";
		ram_buffer(547) := X"1040FFFC";
		ram_buffer(548) := X"00000000";
		ram_buffer(549) := X"AC650008";
		ram_buffer(550) := X"03E00008";
		ram_buffer(551) := X"00000000";
		ram_buffer(552) := X"27BDFFE8";
		ram_buffer(553) := X"AFBF0014";
		ram_buffer(554) := X"0C400AC4";
		ram_buffer(555) := X"00000000";
		ram_buffer(556) := X"10400002";
		ram_buffer(557) := X"24020001";
		ram_buffer(558) := X"AF828054";
		ram_buffer(559) := X"8FBF0014";
		ram_buffer(560) := X"8F82808C";
		ram_buffer(561) := X"24030007";
		ram_buffer(562) := X"AC430000";
		ram_buffer(563) := X"03E00008";
		ram_buffer(564) := X"27BD0018";
		ram_buffer(565) := X"8F828094";
		ram_buffer(566) := X"3C040100";
		ram_buffer(567) := X"8C420004";
		ram_buffer(568) := X"084004DC";
		ram_buffer(569) := X"248454CC";
		ram_buffer(570) := X"03E00008";
		ram_buffer(571) := X"00000000";
		ram_buffer(572) := X"24020001";
		ram_buffer(573) := X"3C030101";
		ram_buffer(574) := X"AF82800C";
		ram_buffer(575) := X"8C625900";
		ram_buffer(576) := X"27BDFFE0";
		ram_buffer(577) := X"8C420004";
		ram_buffer(578) := X"AFB10018";
		ram_buffer(579) := X"3C110101";
		ram_buffer(580) := X"AFB00014";
		ram_buffer(581) := X"AFBF001C";
		ram_buffer(582) := X"00608025";
		ram_buffer(583) := X"26315904";
		ram_buffer(584) := X"2C430008";
		ram_buffer(585) := X"14600014";
		ram_buffer(586) := X"000210C0";
		ram_buffer(587) := X"8F828008";
		ram_buffer(588) := X"00000000";
		ram_buffer(589) := X"10400004";
		ram_buffer(590) := X"00000000";
		ram_buffer(591) := X"AF808008";
		ram_buffer(592) := X"0C40023A";
		ram_buffer(593) := X"00000000";
		ram_buffer(594) := X"AF80800C";
		ram_buffer(595) := X"8F828054";
		ram_buffer(596) := X"00000000";
		ram_buffer(597) := X"10400012";
		ram_buffer(598) := X"00000000";
		ram_buffer(599) := X"8FBF001C";
		ram_buffer(600) := X"8FB10018";
		ram_buffer(601) := X"8FB00014";
		ram_buffer(602) := X"27BD0020";
		ram_buffer(603) := X"AF808054";
		ram_buffer(604) := X"08400B3F";
		ram_buffer(605) := X"00000000";
		ram_buffer(606) := X"02221021";
		ram_buffer(607) := X"8C430000";
		ram_buffer(608) := X"8C440004";
		ram_buffer(609) := X"0060F809";
		ram_buffer(610) := X"00000000";
		ram_buffer(611) := X"8E025900";
		ram_buffer(612) := X"00000000";
		ram_buffer(613) := X"8C420004";
		ram_buffer(614) := X"1000FFE2";
		ram_buffer(615) := X"2C430008";
		ram_buffer(616) := X"8FBF001C";
		ram_buffer(617) := X"8FB10018";
		ram_buffer(618) := X"8FB00014";
		ram_buffer(619) := X"03E00008";
		ram_buffer(620) := X"27BD0020";
		ram_buffer(621) := X"27BDFFE0";
		ram_buffer(622) := X"8F828090";
		ram_buffer(623) := X"3403FFFF";
		ram_buffer(624) := X"AFB00010";
		ram_buffer(625) := X"3C100100";
		ram_buffer(626) := X"AFB20018";
		ram_buffer(627) := X"AFB10014";
		ram_buffer(628) := X"AFBF001C";
		ram_buffer(629) := X"00808825";
		ram_buffer(630) := X"00A09025";
		ram_buffer(631) := X"AC430008";
		ram_buffer(632) := X"261054D8";
		ram_buffer(633) := X"02403025";
		ram_buffer(634) := X"02202825";
		ram_buffer(635) := X"0C4004DC";
		ram_buffer(636) := X"02002025";
		ram_buffer(637) := X"1000FFFC";
		ram_buffer(638) := X"02403025";
		ram_buffer(639) := X"3C020101";
		ram_buffer(640) := X"8C425900";
		ram_buffer(641) := X"240300FF";
		ram_buffer(642) := X"03E00008";
		ram_buffer(643) := X"AC430000";
		ram_buffer(644) := X"3C020101";
		ram_buffer(645) := X"8C425900";
		ram_buffer(646) := X"00000000";
		ram_buffer(647) := X"03E00008";
		ram_buffer(648) := X"AC400000";
		ram_buffer(649) := X"24020001";
		ram_buffer(650) := X"AF828008";
		ram_buffer(651) := X"08400120";
		ram_buffer(652) := X"00000000";
		ram_buffer(653) := X"27BDFFE8";
		ram_buffer(654) := X"AFB00010";
		ram_buffer(655) := X"00808025";
		ram_buffer(656) := X"AFBF0014";
		ram_buffer(657) := X"0C400046";
		ram_buffer(658) := X"00002025";
		ram_buffer(659) := X"3C0344A0";
		ram_buffer(660) := X"3C020101";
		ram_buffer(661) := X"AC435900";
		ram_buffer(662) := X"3C040101";
		ram_buffer(663) := X"3C030101";
		ram_buffer(664) := X"24635904";
		ram_buffer(665) := X"24845944";
		ram_buffer(666) := X"24630008";
		ram_buffer(667) := X"1464FFFE";
		ram_buffer(668) := X"AC60FFF8";
		ram_buffer(669) := X"3C0344A2";
		ram_buffer(670) := X"AF838090";
		ram_buffer(671) := X"3404C350";
		ram_buffer(672) := X"3C0344A1";
		ram_buffer(673) := X"AF83808C";
		ram_buffer(674) := X"AC640004";
		ram_buffer(675) := X"3C030100";
		ram_buffer(676) := X"24425900";
		ram_buffer(677) := X"246308A0";
		ram_buffer(678) := X"AC430004";
		ram_buffer(679) := X"3C0344A4";
		ram_buffer(680) := X"AF838094";
		ram_buffer(681) := X"3C030100";
		ram_buffer(682) := X"246308D4";
		ram_buffer(683) := X"3C050100";
		ram_buffer(684) := X"AC400008";
		ram_buffer(685) := X"AC43001C";
		ram_buffer(686) := X"AC400020";
		ram_buffer(687) := X"24A50878";
		ram_buffer(688) := X"0C4004D9";
		ram_buffer(689) := X"00002025";
		ram_buffer(690) := X"0200F809";
		ram_buffer(691) := X"00000000";
		ram_buffer(692) := X"8F82808C";
		ram_buffer(693) := X"24030003";
		ram_buffer(694) := X"AC430000";
		ram_buffer(695) := X"8F828090";
		ram_buffer(696) := X"24030001";
		ram_buffer(697) := X"0C400DBB";
		ram_buffer(698) := X"AC430008";
		ram_buffer(699) := X"3C040100";
		ram_buffer(700) := X"240500CF";
		ram_buffer(701) := X"0C40026D";
		ram_buffer(702) := X"248454F8";
		ram_buffer(703) := X"00041080";
		ram_buffer(704) := X"3C040101";
		ram_buffer(705) := X"24845944";
		ram_buffer(706) := X"00822021";
		ram_buffer(707) := X"2402001F";
		ram_buffer(708) := X"00452823";
		ram_buffer(709) := X"24020006";
		ram_buffer(710) := X"14400002";
		ram_buffer(711) := X"00A2001A";
		ram_buffer(712) := X"0007000D";
		ram_buffer(713) := X"27BDFFE0";
		ram_buffer(714) := X"00C01825";
		ram_buffer(715) := X"00003825";
		ram_buffer(716) := X"AFA40014";
		ram_buffer(717) := X"2406012C";
		ram_buffer(718) := X"00602025";
		ram_buffer(719) := X"AFBF001C";
		ram_buffer(720) := X"00002812";
		ram_buffer(721) := X"AFA50010";
		ram_buffer(722) := X"0C400D00";
		ram_buffer(723) := X"00002825";
		ram_buffer(724) := X"24030001";
		ram_buffer(725) := X"10430005";
		ram_buffer(726) := X"00001025";
		ram_buffer(727) := X"3C040100";
		ram_buffer(728) := X"240500DD";
		ram_buffer(729) := X"0C40026D";
		ram_buffer(730) := X"248454F8";
		ram_buffer(731) := X"8FBF001C";
		ram_buffer(732) := X"00000000";
		ram_buffer(733) := X"03E00008";
		ram_buffer(734) := X"27BD0020";
		ram_buffer(735) := X"3C030101";
		ram_buffer(736) := X"00042080";
		ram_buffer(737) := X"24625944";
		ram_buffer(738) := X"8F85800C";
		ram_buffer(739) := X"27BDFFE8";
		ram_buffer(740) := X"00441021";
		ram_buffer(741) := X"8C440000";
		ram_buffer(742) := X"10A0000A";
		ram_buffer(743) := X"AFBF0014";
		ram_buffer(744) := X"0C400A5B";
		ram_buffer(745) := X"00000000";
		ram_buffer(746) := X"10400002";
		ram_buffer(747) := X"24020001";
		ram_buffer(748) := X"AF828054";
		ram_buffer(749) := X"8FBF0014";
		ram_buffer(750) := X"00001025";
		ram_buffer(751) := X"03E00008";
		ram_buffer(752) := X"27BD0018";
		ram_buffer(753) := X"0C400F0C";
		ram_buffer(754) := X"00000000";
		ram_buffer(755) := X"1000FFF9";
		ram_buffer(756) := X"00000000";
		ram_buffer(757) := X"3C020101";
		ram_buffer(758) := X"24425944";
		ram_buffer(759) := X"00042080";
		ram_buffer(760) := X"00822021";
		ram_buffer(761) := X"8C840000";
		ram_buffer(762) := X"27BDFFE8";
		ram_buffer(763) := X"AFBF0014";
		ram_buffer(764) := X"0C400EC5";
		ram_buffer(765) := X"00000000";
		ram_buffer(766) := X"8FBF0014";
		ram_buffer(767) := X"00001025";
		ram_buffer(768) := X"03E00008";
		ram_buffer(769) := X"27BD0018";
		ram_buffer(770) := X"08400120";
		ram_buffer(771) := X"00000000";
		ram_buffer(772) := X"240203E8";
		ram_buffer(773) := X"00820018";
		ram_buffer(774) := X"00002012";
		ram_buffer(775) := X"08400FE4";
		ram_buffer(776) := X"00000000";
		ram_buffer(777) := X"27BDFFE8";
		ram_buffer(778) := X"00003025";
		ram_buffer(779) := X"24050010";
		ram_buffer(780) := X"AFB00010";
		ram_buffer(781) := X"00808025";
		ram_buffer(782) := X"24040001";
		ram_buffer(783) := X"AFBF0014";
		ram_buffer(784) := X"0C40061D";
		ram_buffer(785) := X"00108080";
		ram_buffer(786) := X"27848088";
		ram_buffer(787) := X"00902021";
		ram_buffer(788) := X"14400005";
		ram_buffer(789) := X"AC820000";
		ram_buffer(790) := X"3C040100";
		ram_buffer(791) := X"24050116";
		ram_buffer(792) := X"0C40026D";
		ram_buffer(793) := X"248454F8";
		ram_buffer(794) := X"8FBF0014";
		ram_buffer(795) := X"8FB00010";
		ram_buffer(796) := X"00001025";
		ram_buffer(797) := X"03E00008";
		ram_buffer(798) := X"27BD0018";
		ram_buffer(799) := X"8F82800C";
		ram_buffer(800) := X"27BDFFE0";
		ram_buffer(801) := X"00042080";
		ram_buffer(802) := X"10400013";
		ram_buffer(803) := X"AFBF001C";
		ram_buffer(804) := X"27828088";
		ram_buffer(805) := X"00442021";
		ram_buffer(806) := X"8C840000";
		ram_buffer(807) := X"00003825";
		ram_buffer(808) := X"27A60010";
		ram_buffer(809) := X"0C40073B";
		ram_buffer(810) := X"AFA00010";
		ram_buffer(811) := X"8FA30010";
		ram_buffer(812) := X"00000000";
		ram_buffer(813) := X"10600003";
		ram_buffer(814) := X"24030001";
		ram_buffer(815) := X"AF838054";
		ram_buffer(816) := X"24030001";
		ram_buffer(817) := X"1043000C";
		ram_buffer(818) := X"3C040100";
		ram_buffer(819) := X"2405012A";
		ram_buffer(820) := X"0C40026D";
		ram_buffer(821) := X"248454F8";
		ram_buffer(822) := X"27828088";
		ram_buffer(823) := X"00442021";
		ram_buffer(824) := X"8C840000";
		ram_buffer(825) := X"00003825";
		ram_buffer(826) := X"0C40065F";
		ram_buffer(827) := X"2406FFFF";
		ram_buffer(828) := X"1000FFF4";
		ram_buffer(829) := X"24030001";
		ram_buffer(830) := X"8FBF001C";
		ram_buffer(831) := X"00001025";
		ram_buffer(832) := X"03E00008";
		ram_buffer(833) := X"27BD0020";
		ram_buffer(834) := X"8F82800C";
		ram_buffer(835) := X"27BDFFE0";
		ram_buffer(836) := X"00042080";
		ram_buffer(837) := X"10400012";
		ram_buffer(838) := X"AFBF001C";
		ram_buffer(839) := X"27828088";
		ram_buffer(840) := X"00442021";
		ram_buffer(841) := X"8C840000";
		ram_buffer(842) := X"27A60010";
		ram_buffer(843) := X"0C4008AE";
		ram_buffer(844) := X"AFA00010";
		ram_buffer(845) := X"8FA30010";
		ram_buffer(846) := X"00000000";
		ram_buffer(847) := X"10600003";
		ram_buffer(848) := X"24030001";
		ram_buffer(849) := X"AF838054";
		ram_buffer(850) := X"24030001";
		ram_buffer(851) := X"1043000C";
		ram_buffer(852) := X"3C040100";
		ram_buffer(853) := X"2405013E";
		ram_buffer(854) := X"0C40026D";
		ram_buffer(855) := X"248454F8";
		ram_buffer(856) := X"27828088";
		ram_buffer(857) := X"00442021";
		ram_buffer(858) := X"8C840000";
		ram_buffer(859) := X"00003825";
		ram_buffer(860) := X"0C4007D5";
		ram_buffer(861) := X"2406FFFF";
		ram_buffer(862) := X"1000FFF4";
		ram_buffer(863) := X"24030001";
		ram_buffer(864) := X"8FBF001C";
		ram_buffer(865) := X"00001025";
		ram_buffer(866) := X"03E00008";
		ram_buffer(867) := X"27BD0020";
		ram_buffer(868) := X"27BDFFE8";
		ram_buffer(869) := X"24050001";
		ram_buffer(870) := X"AFB00010";
		ram_buffer(871) := X"00808025";
		ram_buffer(872) := X"24040001";
		ram_buffer(873) := X"AFBF0014";
		ram_buffer(874) := X"0C400641";
		ram_buffer(875) := X"00108080";
		ram_buffer(876) := X"2784809C";
		ram_buffer(877) := X"00902021";
		ram_buffer(878) := X"14400005";
		ram_buffer(879) := X"AC820000";
		ram_buffer(880) := X"3C040100";
		ram_buffer(881) := X"2405014A";
		ram_buffer(882) := X"0C40026D";
		ram_buffer(883) := X"248454F8";
		ram_buffer(884) := X"8FBF0014";
		ram_buffer(885) := X"8FB00010";
		ram_buffer(886) := X"00001025";
		ram_buffer(887) := X"03E00008";
		ram_buffer(888) := X"27BD0018";
		ram_buffer(889) := X"8F82800C";
		ram_buffer(890) := X"27BDFFE0";
		ram_buffer(891) := X"00042080";
		ram_buffer(892) := X"10400013";
		ram_buffer(893) := X"AFBF001C";
		ram_buffer(894) := X"2782809C";
		ram_buffer(895) := X"00442021";
		ram_buffer(896) := X"8C840000";
		ram_buffer(897) := X"27A60010";
		ram_buffer(898) := X"00002825";
		ram_buffer(899) := X"0C4008AE";
		ram_buffer(900) := X"AFA00010";
		ram_buffer(901) := X"8FA30010";
		ram_buffer(902) := X"00000000";
		ram_buffer(903) := X"10600003";
		ram_buffer(904) := X"24030001";
		ram_buffer(905) := X"AF838054";
		ram_buffer(906) := X"24030001";
		ram_buffer(907) := X"1043000D";
		ram_buffer(908) := X"3C040100";
		ram_buffer(909) := X"2405015E";
		ram_buffer(910) := X"0C40026D";
		ram_buffer(911) := X"248454F8";
		ram_buffer(912) := X"2782809C";
		ram_buffer(913) := X"00442021";
		ram_buffer(914) := X"8C840000";
		ram_buffer(915) := X"00003825";
		ram_buffer(916) := X"2406FFFF";
		ram_buffer(917) := X"0C4007D5";
		ram_buffer(918) := X"00002825";
		ram_buffer(919) := X"1000FFF3";
		ram_buffer(920) := X"24030001";
		ram_buffer(921) := X"8FBF001C";
		ram_buffer(922) := X"00001025";
		ram_buffer(923) := X"03E00008";
		ram_buffer(924) := X"27BD0020";
		ram_buffer(925) := X"8F82800C";
		ram_buffer(926) := X"27BDFFE0";
		ram_buffer(927) := X"00042080";
		ram_buffer(928) := X"10400012";
		ram_buffer(929) := X"AFBF001C";
		ram_buffer(930) := X"2782809C";
		ram_buffer(931) := X"00442021";
		ram_buffer(932) := X"8C840000";
		ram_buffer(933) := X"27A50010";
		ram_buffer(934) := X"0C400791";
		ram_buffer(935) := X"AFA00010";
		ram_buffer(936) := X"8FA30010";
		ram_buffer(937) := X"00000000";
		ram_buffer(938) := X"10600003";
		ram_buffer(939) := X"24030001";
		ram_buffer(940) := X"AF838054";
		ram_buffer(941) := X"24030001";
		ram_buffer(942) := X"1043000D";
		ram_buffer(943) := X"3C040100";
		ram_buffer(944) := X"24050172";
		ram_buffer(945) := X"0C40026D";
		ram_buffer(946) := X"248454F8";
		ram_buffer(947) := X"2782809C";
		ram_buffer(948) := X"00442021";
		ram_buffer(949) := X"8C840000";
		ram_buffer(950) := X"00003825";
		ram_buffer(951) := X"00003025";
		ram_buffer(952) := X"0C40065F";
		ram_buffer(953) := X"00002825";
		ram_buffer(954) := X"1000FFF3";
		ram_buffer(955) := X"24030001";
		ram_buffer(956) := X"8FBF001C";
		ram_buffer(957) := X"00001025";
		ram_buffer(958) := X"03E00008";
		ram_buffer(959) := X"27BD0020";
		ram_buffer(960) := X"03E00008";
		ram_buffer(961) := X"00001025";
		ram_buffer(962) := X"27BDFFE0";
		ram_buffer(963) := X"AFB00014";
		ram_buffer(964) := X"00808025";
		ram_buffer(965) := X"24040080";
		ram_buffer(966) := X"AFB10018";
		ram_buffer(967) := X"AFBF001C";
		ram_buffer(968) := X"00A08825";
		ram_buffer(969) := X"0C4012E8";
		ram_buffer(970) := X"00108080";
		ram_buffer(971) := X"27848098";
		ram_buffer(972) := X"00902021";
		ram_buffer(973) := X"AC820000";
		ram_buffer(974) := X"14400005";
		ram_buffer(975) := X"AE220000";
		ram_buffer(976) := X"3C040100";
		ram_buffer(977) := X"24050189";
		ram_buffer(978) := X"0C40026D";
		ram_buffer(979) := X"248454F8";
		ram_buffer(980) := X"8FBF001C";
		ram_buffer(981) := X"8FB10018";
		ram_buffer(982) := X"8FB00014";
		ram_buffer(983) := X"00001025";
		ram_buffer(984) := X"03E00008";
		ram_buffer(985) := X"27BD0020";
		ram_buffer(986) := X"27828098";
		ram_buffer(987) := X"00042080";
		ram_buffer(988) := X"00442021";
		ram_buffer(989) := X"8C840000";
		ram_buffer(990) := X"27BDFFE8";
		ram_buffer(991) := X"24020001";
		ram_buffer(992) := X"14850004";
		ram_buffer(993) := X"AFBF0014";
		ram_buffer(994) := X"0C40135A";
		ram_buffer(995) := X"00000000";
		ram_buffer(996) := X"00001025";
		ram_buffer(997) := X"8FBF0014";
		ram_buffer(998) := X"00000000";
		ram_buffer(999) := X"03E00008";
		ram_buffer(1000) := X"27BD0018";
		ram_buffer(1001) := X"24020001";
		ram_buffer(1002) := X"14400002";
		ram_buffer(1003) := X"0082001B";
		ram_buffer(1004) := X"0007000D";
		ram_buffer(1005) := X"00001812";
		ram_buffer(1006) := X"0065182B";
		ram_buffer(1007) := X"10600006";
		ram_buffer(1008) := X"00450018";
		ram_buffer(1009) := X"00004025";
		ram_buffer(1010) := X"14400006";
		ram_buffer(1011) := X"00000000";
		ram_buffer(1012) := X"03E00008";
		ram_buffer(1013) := X"A0E00000";
		ram_buffer(1014) := X"00001012";
		ram_buffer(1015) := X"1000FFF2";
		ram_buffer(1016) := X"00000000";
		ram_buffer(1017) := X"14400002";
		ram_buffer(1018) := X"0082001B";
		ram_buffer(1019) := X"0007000D";
		ram_buffer(1020) := X"00002010";
		ram_buffer(1021) := X"00004812";
		ram_buffer(1022) := X"00000000";
		ram_buffer(1023) := X"00000000";
		ram_buffer(1024) := X"14A00002";
		ram_buffer(1025) := X"0045001B";
		ram_buffer(1026) := X"0007000D";
		ram_buffer(1027) := X"00001012";
		ram_buffer(1028) := X"15000005";
		ram_buffer(1029) := X"292A000A";
		ram_buffer(1030) := X"1D200004";
		ram_buffer(1031) := X"24EB0001";
		ram_buffer(1032) := X"1440FFE9";
		ram_buffer(1033) := X"00000000";
		ram_buffer(1034) := X"24EB0001";
		ram_buffer(1035) := X"15400004";
		ram_buffer(1036) := X"24030030";
		ram_buffer(1037) := X"14C00002";
		ram_buffer(1038) := X"24030037";
		ram_buffer(1039) := X"24030057";
		ram_buffer(1040) := X"00691821";
		ram_buffer(1041) := X"A0E30000";
		ram_buffer(1042) := X"25080001";
		ram_buffer(1043) := X"1000FFDE";
		ram_buffer(1044) := X"01603825";
		ram_buffer(1045) := X"27BDFFD8";
		ram_buffer(1046) := X"AFB40020";
		ram_buffer(1047) := X"AFB3001C";
		ram_buffer(1048) := X"AFB20018";
		ram_buffer(1049) := X"AFB10014";
		ram_buffer(1050) := X"AFBF0024";
		ram_buffer(1051) := X"AFB00010";
		ram_buffer(1052) := X"00809025";
		ram_buffer(1053) := X"00A09825";
		ram_buffer(1054) := X"8FB10038";
		ram_buffer(1055) := X"10E00002";
		ram_buffer(1056) := X"24140020";
		ram_buffer(1057) := X"24140030";
		ram_buffer(1058) := X"02201025";
		ram_buffer(1059) := X"24420001";
		ram_buffer(1060) := X"8043FFFF";
		ram_buffer(1061) := X"00000000";
		ram_buffer(1062) := X"14600009";
		ram_buffer(1063) := X"00C08025";
		ram_buffer(1064) := X"1A000009";
		ram_buffer(1065) := X"02802825";
		ram_buffer(1066) := X"0260F809";
		ram_buffer(1067) := X"02402025";
		ram_buffer(1068) := X"1000FFFB";
		ram_buffer(1069) := X"2610FFFF";
		ram_buffer(1070) := X"1000FFF4";
		ram_buffer(1071) := X"24C6FFFF";
		ram_buffer(1072) := X"1CC0FFFD";
		ram_buffer(1073) := X"00000000";
		ram_buffer(1074) := X"26310001";
		ram_buffer(1075) := X"8225FFFF";
		ram_buffer(1076) := X"00000000";
		ram_buffer(1077) := X"14A00009";
		ram_buffer(1078) := X"00000000";
		ram_buffer(1079) := X"8FBF0024";
		ram_buffer(1080) := X"8FB40020";
		ram_buffer(1081) := X"8FB3001C";
		ram_buffer(1082) := X"8FB20018";
		ram_buffer(1083) := X"8FB10014";
		ram_buffer(1084) := X"8FB00010";
		ram_buffer(1085) := X"03E00008";
		ram_buffer(1086) := X"27BD0028";
		ram_buffer(1087) := X"0260F809";
		ram_buffer(1088) := X"02402025";
		ram_buffer(1089) := X"1000FFF1";
		ram_buffer(1090) := X"26310001";
		ram_buffer(1091) := X"8C820000";
		ram_buffer(1092) := X"00000000";
		ram_buffer(1093) := X"24430001";
		ram_buffer(1094) := X"AC830000";
		ram_buffer(1095) := X"03E00008";
		ram_buffer(1096) := X"A0450000";
		ram_buffer(1097) := X"27BDFFB8";
		ram_buffer(1098) := X"AFB5003C";
		ram_buffer(1099) := X"AFB40038";
		ram_buffer(1100) := X"AFB30034";
		ram_buffer(1101) := X"AFB20030";
		ram_buffer(1102) := X"AFB1002C";
		ram_buffer(1103) := X"AFB00028";
		ram_buffer(1104) := X"AFBF0044";
		ram_buffer(1105) := X"AFB60040";
		ram_buffer(1106) := X"00809025";
		ram_buffer(1107) := X"00A09825";
		ram_buffer(1108) := X"00C08825";
		ram_buffer(1109) := X"00E08025";
		ram_buffer(1110) := X"24140025";
		ram_buffer(1111) := X"24150030";
		ram_buffer(1112) := X"82250000";
		ram_buffer(1113) := X"00000000";
		ram_buffer(1114) := X"10A00035";
		ram_buffer(1115) := X"00000000";
		ram_buffer(1116) := X"10B40006";
		ram_buffer(1117) := X"00000000";
		ram_buffer(1118) := X"26310001";
		ram_buffer(1119) := X"0260F809";
		ram_buffer(1120) := X"02402025";
		ram_buffer(1121) := X"1000FFF6";
		ram_buffer(1122) := X"00000000";
		ram_buffer(1123) := X"82260001";
		ram_buffer(1124) := X"00000000";
		ram_buffer(1125) := X"10D50015";
		ram_buffer(1126) := X"240D0001";
		ram_buffer(1127) := X"26310002";
		ram_buffer(1128) := X"00006825";
		ram_buffer(1129) := X"24C2FFD0";
		ram_buffer(1130) := X"304200FF";
		ram_buffer(1131) := X"2C42000A";
		ram_buffer(1132) := X"10400018";
		ram_buffer(1133) := X"00006025";
		ram_buffer(1134) := X"30C200FF";
		ram_buffer(1135) := X"2443FFD0";
		ram_buffer(1136) := X"2C63000A";
		ram_buffer(1137) := X"1060000C";
		ram_buffer(1138) := X"2443FF9F";
		ram_buffer(1139) := X"24C3FFD0";
		ram_buffer(1140) := X"000C1080";
		ram_buffer(1141) := X"004C6021";
		ram_buffer(1142) := X"000C6040";
		ram_buffer(1143) := X"26310001";
		ram_buffer(1144) := X"8226FFFF";
		ram_buffer(1145) := X"1000FFF4";
		ram_buffer(1146) := X"01836021";
		ram_buffer(1147) := X"82260002";
		ram_buffer(1148) := X"1000FFEC";
		ram_buffer(1149) := X"26310003";
		ram_buffer(1150) := X"2C630006";
		ram_buffer(1151) := X"1060001A";
		ram_buffer(1152) := X"2442FFBF";
		ram_buffer(1153) := X"24C3FFA9";
		ram_buffer(1154) := X"2862000B";
		ram_buffer(1155) := X"1440FFF1";
		ram_buffer(1156) := X"000C1080";
		ram_buffer(1157) := X"24020063";
		ram_buffer(1158) := X"10C20045";
		ram_buffer(1159) := X"28C20064";
		ram_buffer(1160) := X"10400016";
		ram_buffer(1161) := X"24020073";
		ram_buffer(1162) := X"10D4004C";
		ram_buffer(1163) := X"24020058";
		ram_buffer(1164) := X"10C20033";
		ram_buffer(1165) := X"00000000";
		ram_buffer(1166) := X"14C0FFC9";
		ram_buffer(1167) := X"00000000";
		ram_buffer(1168) := X"8FBF0044";
		ram_buffer(1169) := X"8FB60040";
		ram_buffer(1170) := X"8FB5003C";
		ram_buffer(1171) := X"8FB40038";
		ram_buffer(1172) := X"8FB30034";
		ram_buffer(1173) := X"8FB20030";
		ram_buffer(1174) := X"8FB1002C";
		ram_buffer(1175) := X"8FB00028";
		ram_buffer(1176) := X"03E00008";
		ram_buffer(1177) := X"27BD0048";
		ram_buffer(1178) := X"2C420006";
		ram_buffer(1179) := X"1040FFEA";
		ram_buffer(1180) := X"24020063";
		ram_buffer(1181) := X"1000FFE4";
		ram_buffer(1182) := X"24C3FFC9";
		ram_buffer(1183) := X"10C20032";
		ram_buffer(1184) := X"28C20074";
		ram_buffer(1185) := X"10400019";
		ram_buffer(1186) := X"24020075";
		ram_buffer(1187) := X"24020064";
		ram_buffer(1188) := X"14C2FFB3";
		ram_buffer(1189) := X"26160004";
		ram_buffer(1190) := X"8E040000";
		ram_buffer(1191) := X"00000000";
		ram_buffer(1192) := X"04810005";
		ram_buffer(1193) := X"27A70018";
		ram_buffer(1194) := X"2402002D";
		ram_buffer(1195) := X"00042023";
		ram_buffer(1196) := X"A3A20018";
		ram_buffer(1197) := X"27A70019";
		ram_buffer(1198) := X"00003025";
		ram_buffer(1199) := X"2405000A";
		ram_buffer(1200) := X"0C4003E9";
		ram_buffer(1201) := X"00000000";
		ram_buffer(1202) := X"27A20018";
		ram_buffer(1203) := X"AFA20010";
		ram_buffer(1204) := X"01A03825";
		ram_buffer(1205) := X"01803025";
		ram_buffer(1206) := X"02602825";
		ram_buffer(1207) := X"0C400415";
		ram_buffer(1208) := X"02402025";
		ram_buffer(1209) := X"1000FF9E";
		ram_buffer(1210) := X"02C08025";
		ram_buffer(1211) := X"10C2000A";
		ram_buffer(1212) := X"26160004";
		ram_buffer(1213) := X"24020078";
		ram_buffer(1214) := X"14C2FF99";
		ram_buffer(1215) := X"00000000";
		ram_buffer(1216) := X"38C60058";
		ram_buffer(1217) := X"26160004";
		ram_buffer(1218) := X"27A70018";
		ram_buffer(1219) := X"2CC60001";
		ram_buffer(1220) := X"10000004";
		ram_buffer(1221) := X"24050010";
		ram_buffer(1222) := X"27A70018";
		ram_buffer(1223) := X"00003025";
		ram_buffer(1224) := X"2405000A";
		ram_buffer(1225) := X"8E040000";
		ram_buffer(1226) := X"1000FFE5";
		ram_buffer(1227) := X"00000000";
		ram_buffer(1228) := X"82050003";
		ram_buffer(1229) := X"02402025";
		ram_buffer(1230) := X"0260F809";
		ram_buffer(1231) := X"26160004";
		ram_buffer(1232) := X"1000FF87";
		ram_buffer(1233) := X"02C08025";
		ram_buffer(1234) := X"8E020000";
		ram_buffer(1235) := X"26160004";
		ram_buffer(1236) := X"AFA20010";
		ram_buffer(1237) := X"1000FFDF";
		ram_buffer(1238) := X"00003825";
		ram_buffer(1239) := X"1000FF87";
		ram_buffer(1240) := X"24050025";
		ram_buffer(1241) := X"AF858014";
		ram_buffer(1242) := X"03E00008";
		ram_buffer(1243) := X"AF848010";
		ram_buffer(1244) := X"27BDFFE0";
		ram_buffer(1245) := X"AFA50024";
		ram_buffer(1246) := X"AFA60028";
		ram_buffer(1247) := X"8F858014";
		ram_buffer(1248) := X"00803025";
		ram_buffer(1249) := X"8F848010";
		ram_buffer(1250) := X"AFA7002C";
		ram_buffer(1251) := X"27A70024";
		ram_buffer(1252) := X"AFBF001C";
		ram_buffer(1253) := X"0C400449";
		ram_buffer(1254) := X"AFA70010";
		ram_buffer(1255) := X"8FBF001C";
		ram_buffer(1256) := X"00000000";
		ram_buffer(1257) := X"03E00008";
		ram_buffer(1258) := X"27BD0020";
		ram_buffer(1259) := X"27BDFFE0";
		ram_buffer(1260) := X"AFA60028";
		ram_buffer(1261) := X"00A03025";
		ram_buffer(1262) := X"3C050100";
		ram_buffer(1263) := X"AFA40020";
		ram_buffer(1264) := X"AFA7002C";
		ram_buffer(1265) := X"27A40020";
		ram_buffer(1266) := X"27A70028";
		ram_buffer(1267) := X"24A5110C";
		ram_buffer(1268) := X"AFBF001C";
		ram_buffer(1269) := X"0C400449";
		ram_buffer(1270) := X"AFA70010";
		ram_buffer(1271) := X"8FA20020";
		ram_buffer(1272) := X"00000000";
		ram_buffer(1273) := X"A0400000";
		ram_buffer(1274) := X"8FBF001C";
		ram_buffer(1275) := X"00000000";
		ram_buffer(1276) := X"03E00008";
		ram_buffer(1277) := X"27BD0020";
		ram_buffer(1278) := X"10C0000D";
		ram_buffer(1279) := X"00C53021";
		ram_buffer(1280) := X"2402FFF0";
		ram_buffer(1281) := X"00C21824";
		ram_buffer(1282) := X"0066302B";
		ram_buffer(1283) := X"00A22824";
		ram_buffer(1284) := X"00063100";
		ram_buffer(1285) := X"24620010";
		ram_buffer(1286) := X"00463021";
		ram_buffer(1287) := X"3C022000";
		ram_buffer(1288) := X"00822021";
		ram_buffer(1289) := X"2402FFF0";
		ram_buffer(1290) := X"14C50003";
		ram_buffer(1291) := X"00A21824";
		ram_buffer(1292) := X"03E00008";
		ram_buffer(1293) := X"00000000";
		ram_buffer(1294) := X"AC830000";
		ram_buffer(1295) := X"AC600000";
		ram_buffer(1296) := X"1000FFF9";
		ram_buffer(1297) := X"24A50010";
		ram_buffer(1298) := X"24820008";
		ram_buffer(1299) := X"2403FFFF";
		ram_buffer(1300) := X"AC820004";
		ram_buffer(1301) := X"AC830008";
		ram_buffer(1302) := X"AC82000C";
		ram_buffer(1303) := X"AC820010";
		ram_buffer(1304) := X"03E00008";
		ram_buffer(1305) := X"AC800000";
		ram_buffer(1306) := X"03E00008";
		ram_buffer(1307) := X"AC800010";
		ram_buffer(1308) := X"8C820004";
		ram_buffer(1309) := X"00000000";
		ram_buffer(1310) := X"8C430008";
		ram_buffer(1311) := X"ACA20004";
		ram_buffer(1312) := X"ACA30008";
		ram_buffer(1313) := X"8C430008";
		ram_buffer(1314) := X"00000000";
		ram_buffer(1315) := X"AC650004";
		ram_buffer(1316) := X"AC450008";
		ram_buffer(1317) := X"8C820000";
		ram_buffer(1318) := X"ACA40010";
		ram_buffer(1319) := X"24420001";
		ram_buffer(1320) := X"03E00008";
		ram_buffer(1321) := X"AC820000";
		ram_buffer(1322) := X"8CA60000";
		ram_buffer(1323) := X"2403FFFF";
		ram_buffer(1324) := X"14C3000F";
		ram_buffer(1325) := X"24820008";
		ram_buffer(1326) := X"8C820010";
		ram_buffer(1327) := X"00000000";
		ram_buffer(1328) := X"8C430004";
		ram_buffer(1329) := X"00000000";
		ram_buffer(1330) := X"ACA30004";
		ram_buffer(1331) := X"AC650008";
		ram_buffer(1332) := X"ACA20008";
		ram_buffer(1333) := X"AC450004";
		ram_buffer(1334) := X"8C820000";
		ram_buffer(1335) := X"ACA40010";
		ram_buffer(1336) := X"24420001";
		ram_buffer(1337) := X"03E00008";
		ram_buffer(1338) := X"AC820000";
		ram_buffer(1339) := X"00E01025";
		ram_buffer(1340) := X"8C470004";
		ram_buffer(1341) := X"00000000";
		ram_buffer(1342) := X"8CE30000";
		ram_buffer(1343) := X"00000000";
		ram_buffer(1344) := X"00C3182B";
		ram_buffer(1345) := X"1060FFF9";
		ram_buffer(1346) := X"00000000";
		ram_buffer(1347) := X"1000FFEC";
		ram_buffer(1348) := X"00000000";
		ram_buffer(1349) := X"8C850004";
		ram_buffer(1350) := X"8C820008";
		ram_buffer(1351) := X"8C830010";
		ram_buffer(1352) := X"ACA20008";
		ram_buffer(1353) := X"8C820008";
		ram_buffer(1354) := X"00000000";
		ram_buffer(1355) := X"AC450004";
		ram_buffer(1356) := X"8C650004";
		ram_buffer(1357) := X"00000000";
		ram_buffer(1358) := X"14850002";
		ram_buffer(1359) := X"00000000";
		ram_buffer(1360) := X"AC620004";
		ram_buffer(1361) := X"8C620000";
		ram_buffer(1362) := X"AC800010";
		ram_buffer(1363) := X"2442FFFF";
		ram_buffer(1364) := X"03E00008";
		ram_buffer(1365) := X"AC620000";
		ram_buffer(1366) := X"27BDFFE0";
		ram_buffer(1367) := X"AFB20018";
		ram_buffer(1368) := X"00C09025";
		ram_buffer(1369) := X"8C860040";
		ram_buffer(1370) := X"AFB10014";
		ram_buffer(1371) := X"AFB00010";
		ram_buffer(1372) := X"AFBF001C";
		ram_buffer(1373) := X"00808025";
		ram_buffer(1374) := X"8C910038";
		ram_buffer(1375) := X"14C00011";
		ram_buffer(1376) := X"00000000";
		ram_buffer(1377) := X"8C830000";
		ram_buffer(1378) := X"00000000";
		ram_buffer(1379) := X"14600005";
		ram_buffer(1380) := X"00001025";
		ram_buffer(1381) := X"8C840004";
		ram_buffer(1382) := X"0C400C98";
		ram_buffer(1383) := X"00000000";
		ram_buffer(1384) := X"AE000004";
		ram_buffer(1385) := X"8FBF001C";
		ram_buffer(1386) := X"26310001";
		ram_buffer(1387) := X"AE110038";
		ram_buffer(1388) := X"8FB20018";
		ram_buffer(1389) := X"8FB10014";
		ram_buffer(1390) := X"8FB00010";
		ram_buffer(1391) := X"03E00008";
		ram_buffer(1392) := X"27BD0020";
		ram_buffer(1393) := X"16400010";
		ram_buffer(1394) := X"00000000";
		ram_buffer(1395) := X"8C840008";
		ram_buffer(1396) := X"0C401393";
		ram_buffer(1397) := X"00000000";
		ram_buffer(1398) := X"8E020008";
		ram_buffer(1399) := X"8E030040";
		ram_buffer(1400) := X"00000000";
		ram_buffer(1401) := X"00431021";
		ram_buffer(1402) := X"8E030004";
		ram_buffer(1403) := X"AE020008";
		ram_buffer(1404) := X"0043182B";
		ram_buffer(1405) := X"1460FFEB";
		ram_buffer(1406) := X"00001025";
		ram_buffer(1407) := X"8E030000";
		ram_buffer(1408) := X"1000FFE8";
		ram_buffer(1409) := X"AE030008";
		ram_buffer(1410) := X"8C84000C";
		ram_buffer(1411) := X"0C401393";
		ram_buffer(1412) := X"00000000";
		ram_buffer(1413) := X"8E030040";
		ram_buffer(1414) := X"8E02000C";
		ram_buffer(1415) := X"00031823";
		ram_buffer(1416) := X"8E040000";
		ram_buffer(1417) := X"00431021";
		ram_buffer(1418) := X"AE02000C";
		ram_buffer(1419) := X"0044102B";
		ram_buffer(1420) := X"10400005";
		ram_buffer(1421) := X"00000000";
		ram_buffer(1422) := X"8E020004";
		ram_buffer(1423) := X"00000000";
		ram_buffer(1424) := X"00431821";
		ram_buffer(1425) := X"AE03000C";
		ram_buffer(1426) := X"24030002";
		ram_buffer(1427) := X"1643FFD5";
		ram_buffer(1428) := X"00001025";
		ram_buffer(1429) := X"0011182B";
		ram_buffer(1430) := X"1000FFD2";
		ram_buffer(1431) := X"02238823";
		ram_buffer(1432) := X"00801025";
		ram_buffer(1433) := X"8C460040";
		ram_buffer(1434) := X"00000000";
		ram_buffer(1435) := X"10C0000E";
		ram_buffer(1436) := X"00A02025";
		ram_buffer(1437) := X"8C43000C";
		ram_buffer(1438) := X"8C450004";
		ram_buffer(1439) := X"00661821";
		ram_buffer(1440) := X"AC43000C";
		ram_buffer(1441) := X"0065182B";
		ram_buffer(1442) := X"14600004";
		ram_buffer(1443) := X"00000000";
		ram_buffer(1444) := X"8C430000";
		ram_buffer(1445) := X"00000000";
		ram_buffer(1446) := X"AC43000C";
		ram_buffer(1447) := X"8C45000C";
		ram_buffer(1448) := X"08401393";
		ram_buffer(1449) := X"00000000";
		ram_buffer(1450) := X"03E00008";
		ram_buffer(1451) := X"00000000";
		ram_buffer(1452) := X"27BDFFE0";
		ram_buffer(1453) := X"AFB00010";
		ram_buffer(1454) := X"AFB20018";
		ram_buffer(1455) := X"AFB10014";
		ram_buffer(1456) := X"AFBF001C";
		ram_buffer(1457) := X"0C400CD3";
		ram_buffer(1458) := X"00808025";
		ram_buffer(1459) := X"92110045";
		ram_buffer(1460) := X"26120024";
		ram_buffer(1461) := X"00118E00";
		ram_buffer(1462) := X"00118E03";
		ram_buffer(1463) := X"1E200013";
		ram_buffer(1464) := X"2402FFFF";
		ram_buffer(1465) := X"A2020045";
		ram_buffer(1466) := X"0C400CE6";
		ram_buffer(1467) := X"00000000";
		ram_buffer(1468) := X"0C400CD3";
		ram_buffer(1469) := X"00000000";
		ram_buffer(1470) := X"92110044";
		ram_buffer(1471) := X"26120010";
		ram_buffer(1472) := X"00118E00";
		ram_buffer(1473) := X"00118E03";
		ram_buffer(1474) := X"1E200016";
		ram_buffer(1475) := X"2402FFFF";
		ram_buffer(1476) := X"8FBF001C";
		ram_buffer(1477) := X"8FB20018";
		ram_buffer(1478) := X"8FB10014";
		ram_buffer(1479) := X"A2020044";
		ram_buffer(1480) := X"8FB00010";
		ram_buffer(1481) := X"08400CE6";
		ram_buffer(1482) := X"27BD0020";
		ram_buffer(1483) := X"8E020024";
		ram_buffer(1484) := X"00000000";
		ram_buffer(1485) := X"1040FFEB";
		ram_buffer(1486) := X"2402FFFF";
		ram_buffer(1487) := X"0C400BB6";
		ram_buffer(1488) := X"02402025";
		ram_buffer(1489) := X"10400003";
		ram_buffer(1490) := X"00000000";
		ram_buffer(1491) := X"0C400C36";
		ram_buffer(1492) := X"00000000";
		ram_buffer(1493) := X"2631FFFF";
		ram_buffer(1494) := X"00118E00";
		ram_buffer(1495) := X"1000FFDF";
		ram_buffer(1496) := X"00118E03";
		ram_buffer(1497) := X"8E020010";
		ram_buffer(1498) := X"00000000";
		ram_buffer(1499) := X"1040FFE8";
		ram_buffer(1500) := X"2402FFFF";
		ram_buffer(1501) := X"0C400BB6";
		ram_buffer(1502) := X"02402025";
		ram_buffer(1503) := X"10400003";
		ram_buffer(1504) := X"00000000";
		ram_buffer(1505) := X"0C400C36";
		ram_buffer(1506) := X"00000000";
		ram_buffer(1507) := X"2631FFFF";
		ram_buffer(1508) := X"00118E00";
		ram_buffer(1509) := X"1000FFDC";
		ram_buffer(1510) := X"00118E03";
		ram_buffer(1511) := X"27BDFFE0";
		ram_buffer(1512) := X"AFB10018";
		ram_buffer(1513) := X"AFB00014";
		ram_buffer(1514) := X"AFBF001C";
		ram_buffer(1515) := X"00808025";
		ram_buffer(1516) := X"14800005";
		ram_buffer(1517) := X"00A08825";
		ram_buffer(1518) := X"3C040100";
		ram_buffer(1519) := X"2405011B";
		ram_buffer(1520) := X"0C40026D";
		ram_buffer(1521) := X"24845514";
		ram_buffer(1522) := X"0C400CD3";
		ram_buffer(1523) := X"00000000";
		ram_buffer(1524) := X"8E050040";
		ram_buffer(1525) := X"8E03003C";
		ram_buffer(1526) := X"8E040000";
		ram_buffer(1527) := X"00A30018";
		ram_buffer(1528) := X"AE000038";
		ram_buffer(1529) := X"AE040008";
		ram_buffer(1530) := X"00001012";
		ram_buffer(1531) := X"00821821";
		ram_buffer(1532) := X"00451023";
		ram_buffer(1533) := X"00821021";
		ram_buffer(1534) := X"AE02000C";
		ram_buffer(1535) := X"2402FFFF";
		ram_buffer(1536) := X"A2020044";
		ram_buffer(1537) := X"AE030004";
		ram_buffer(1538) := X"A2020045";
		ram_buffer(1539) := X"16200013";
		ram_buffer(1540) := X"00000000";
		ram_buffer(1541) := X"8E020010";
		ram_buffer(1542) := X"00000000";
		ram_buffer(1543) := X"10400007";
		ram_buffer(1544) := X"00000000";
		ram_buffer(1545) := X"0C400BB6";
		ram_buffer(1546) := X"26040010";
		ram_buffer(1547) := X"10400003";
		ram_buffer(1548) := X"00000000";
		ram_buffer(1549) := X"0C400120";
		ram_buffer(1550) := X"00000000";
		ram_buffer(1551) := X"0C400CE6";
		ram_buffer(1552) := X"00000000";
		ram_buffer(1553) := X"8FBF001C";
		ram_buffer(1554) := X"8FB10018";
		ram_buffer(1555) := X"8FB00014";
		ram_buffer(1556) := X"24020001";
		ram_buffer(1557) := X"03E00008";
		ram_buffer(1558) := X"27BD0020";
		ram_buffer(1559) := X"0C400512";
		ram_buffer(1560) := X"26040010";
		ram_buffer(1561) := X"0C400512";
		ram_buffer(1562) := X"26040024";
		ram_buffer(1563) := X"1000FFF3";
		ram_buffer(1564) := X"00000000";
		ram_buffer(1565) := X"27BDFFE0";
		ram_buffer(1566) := X"AFB20018";
		ram_buffer(1567) := X"AFB10014";
		ram_buffer(1568) := X"AFBF001C";
		ram_buffer(1569) := X"AFB00010";
		ram_buffer(1570) := X"00809025";
		ram_buffer(1571) := X"14800005";
		ram_buffer(1572) := X"00A08825";
		ram_buffer(1573) := X"3C040100";
		ram_buffer(1574) := X"24050188";
		ram_buffer(1575) := X"0C40026D";
		ram_buffer(1576) := X"24845514";
		ram_buffer(1577) := X"02510018";
		ram_buffer(1578) := X"00002012";
		ram_buffer(1579) := X"0C4012E8";
		ram_buffer(1580) := X"24840048";
		ram_buffer(1581) := X"10400009";
		ram_buffer(1582) := X"00408025";
		ram_buffer(1583) := X"1620000E";
		ram_buffer(1584) := X"00000000";
		ram_buffer(1585) := X"AE020000";
		ram_buffer(1586) := X"AE12003C";
		ram_buffer(1587) := X"AE110040";
		ram_buffer(1588) := X"24050001";
		ram_buffer(1589) := X"0C4005E7";
		ram_buffer(1590) := X"02002025";
		ram_buffer(1591) := X"8FBF001C";
		ram_buffer(1592) := X"02001025";
		ram_buffer(1593) := X"8FB20018";
		ram_buffer(1594) := X"8FB10014";
		ram_buffer(1595) := X"8FB00010";
		ram_buffer(1596) := X"03E00008";
		ram_buffer(1597) := X"27BD0020";
		ram_buffer(1598) := X"24420048";
		ram_buffer(1599) := X"1000FFF2";
		ram_buffer(1600) := X"AE020000";
		ram_buffer(1601) := X"27BDFFE0";
		ram_buffer(1602) := X"AFB10018";
		ram_buffer(1603) := X"AFB00014";
		ram_buffer(1604) := X"AFBF001C";
		ram_buffer(1605) := X"00808025";
		ram_buffer(1606) := X"14800005";
		ram_buffer(1607) := X"00A08825";
		ram_buffer(1608) := X"3C040100";
		ram_buffer(1609) := X"240502BD";
		ram_buffer(1610) := X"0C40026D";
		ram_buffer(1611) := X"24845514";
		ram_buffer(1612) := X"0211102B";
		ram_buffer(1613) := X"10400006";
		ram_buffer(1614) := X"24060002";
		ram_buffer(1615) := X"3C040100";
		ram_buffer(1616) := X"240502BE";
		ram_buffer(1617) := X"0C40026D";
		ram_buffer(1618) := X"24845514";
		ram_buffer(1619) := X"24060002";
		ram_buffer(1620) := X"00002825";
		ram_buffer(1621) := X"0C40061D";
		ram_buffer(1622) := X"02002025";
		ram_buffer(1623) := X"10400002";
		ram_buffer(1624) := X"00000000";
		ram_buffer(1625) := X"AC510038";
		ram_buffer(1626) := X"8FBF001C";
		ram_buffer(1627) := X"8FB10018";
		ram_buffer(1628) := X"8FB00014";
		ram_buffer(1629) := X"03E00008";
		ram_buffer(1630) := X"27BD0020";
		ram_buffer(1631) := X"27BDFFC0";
		ram_buffer(1632) := X"AFB30028";
		ram_buffer(1633) := X"AFB10020";
		ram_buffer(1634) := X"AFB0001C";
		ram_buffer(1635) := X"AFBF003C";
		ram_buffer(1636) := X"AFB70038";
		ram_buffer(1637) := X"AFB60034";
		ram_buffer(1638) := X"AFB50030";
		ram_buffer(1639) := X"AFB4002C";
		ram_buffer(1640) := X"AFB20024";
		ram_buffer(1641) := X"00808025";
		ram_buffer(1642) := X"00A09825";
		ram_buffer(1643) := X"AFA60048";
		ram_buffer(1644) := X"14800005";
		ram_buffer(1645) := X"00E08825";
		ram_buffer(1646) := X"3C040100";
		ram_buffer(1647) := X"240502D9";
		ram_buffer(1648) := X"0C40026D";
		ram_buffer(1649) := X"24845514";
		ram_buffer(1650) := X"16600006";
		ram_buffer(1651) := X"24020002";
		ram_buffer(1652) := X"8E020040";
		ram_buffer(1653) := X"00000000";
		ram_buffer(1654) := X"14400083";
		ram_buffer(1655) := X"240502DA";
		ram_buffer(1656) := X"24020002";
		ram_buffer(1657) := X"16220005";
		ram_buffer(1658) := X"24020001";
		ram_buffer(1659) := X"8E03003C";
		ram_buffer(1660) := X"00000000";
		ram_buffer(1661) := X"14620081";
		ram_buffer(1662) := X"3C040100";
		ram_buffer(1663) := X"0C400C4D";
		ram_buffer(1664) := X"00000000";
		ram_buffer(1665) := X"14400009";
		ram_buffer(1666) := X"0000B025";
		ram_buffer(1667) := X"8FA20048";
		ram_buffer(1668) := X"00000000";
		ram_buffer(1669) := X"10400005";
		ram_buffer(1670) := X"3C040100";
		ram_buffer(1671) := X"240502DE";
		ram_buffer(1672) := X"0C40026D";
		ram_buffer(1673) := X"24845514";
		ram_buffer(1674) := X"0000B025";
		ram_buffer(1675) := X"24150002";
		ram_buffer(1676) := X"2412FFFF";
		ram_buffer(1677) := X"1000003B";
		ram_buffer(1678) := X"26140010";
		ram_buffer(1679) := X"8FA20048";
		ram_buffer(1680) := X"00000000";
		ram_buffer(1681) := X"14400005";
		ram_buffer(1682) := X"00000000";
		ram_buffer(1683) := X"0C400CE6";
		ram_buffer(1684) := X"00000000";
		ram_buffer(1685) := X"1000004D";
		ram_buffer(1686) := X"00001025";
		ram_buffer(1687) := X"16C00003";
		ram_buffer(1688) := X"00000000";
		ram_buffer(1689) := X"0C400C24";
		ram_buffer(1690) := X"27A40010";
		ram_buffer(1691) := X"0C400CE6";
		ram_buffer(1692) := X"00000000";
		ram_buffer(1693) := X"0C400A98";
		ram_buffer(1694) := X"00000000";
		ram_buffer(1695) := X"0C400CD3";
		ram_buffer(1696) := X"00000000";
		ram_buffer(1697) := X"92020044";
		ram_buffer(1698) := X"00000000";
		ram_buffer(1699) := X"00021600";
		ram_buffer(1700) := X"00021603";
		ram_buffer(1701) := X"14520002";
		ram_buffer(1702) := X"00000000";
		ram_buffer(1703) := X"A2000044";
		ram_buffer(1704) := X"92020045";
		ram_buffer(1705) := X"00000000";
		ram_buffer(1706) := X"00021600";
		ram_buffer(1707) := X"00021603";
		ram_buffer(1708) := X"14520002";
		ram_buffer(1709) := X"00000000";
		ram_buffer(1710) := X"A2000045";
		ram_buffer(1711) := X"0C400CE6";
		ram_buffer(1712) := X"00000000";
		ram_buffer(1713) := X"27A50048";
		ram_buffer(1714) := X"0C4010AC";
		ram_buffer(1715) := X"27A40010";
		ram_buffer(1716) := X"1440003F";
		ram_buffer(1717) := X"00000000";
		ram_buffer(1718) := X"0C400CD3";
		ram_buffer(1719) := X"00000000";
		ram_buffer(1720) := X"8E170038";
		ram_buffer(1721) := X"8E16003C";
		ram_buffer(1722) := X"0C400CE6";
		ram_buffer(1723) := X"00000000";
		ram_buffer(1724) := X"16F60031";
		ram_buffer(1725) := X"00000000";
		ram_buffer(1726) := X"8FA50048";
		ram_buffer(1727) := X"0C400B7C";
		ram_buffer(1728) := X"02802025";
		ram_buffer(1729) := X"0C4005AC";
		ram_buffer(1730) := X"02002025";
		ram_buffer(1731) := X"0C400F41";
		ram_buffer(1732) := X"00000000";
		ram_buffer(1733) := X"14400003";
		ram_buffer(1734) := X"24160001";
		ram_buffer(1735) := X"0C400120";
		ram_buffer(1736) := X"00000000";
		ram_buffer(1737) := X"0C400CD3";
		ram_buffer(1738) := X"00000000";
		ram_buffer(1739) := X"8E020038";
		ram_buffer(1740) := X"8E03003C";
		ram_buffer(1741) := X"00000000";
		ram_buffer(1742) := X"0043102B";
		ram_buffer(1743) := X"14400003";
		ram_buffer(1744) := X"02203025";
		ram_buffer(1745) := X"1635FFBD";
		ram_buffer(1746) := X"00000000";
		ram_buffer(1747) := X"02602825";
		ram_buffer(1748) := X"0C400556";
		ram_buffer(1749) := X"02002025";
		ram_buffer(1750) := X"8E030024";
		ram_buffer(1751) := X"00000000";
		ram_buffer(1752) := X"10600003";
		ram_buffer(1753) := X"00000000";
		ram_buffer(1754) := X"0C400BB6";
		ram_buffer(1755) := X"26040024";
		ram_buffer(1756) := X"10400003";
		ram_buffer(1757) := X"00000000";
		ram_buffer(1758) := X"0C400120";
		ram_buffer(1759) := X"00000000";
		ram_buffer(1760) := X"0C400CE6";
		ram_buffer(1761) := X"00000000";
		ram_buffer(1762) := X"24020001";
		ram_buffer(1763) := X"8FBF003C";
		ram_buffer(1764) := X"8FB70038";
		ram_buffer(1765) := X"8FB60034";
		ram_buffer(1766) := X"8FB50030";
		ram_buffer(1767) := X"8FB4002C";
		ram_buffer(1768) := X"8FB30028";
		ram_buffer(1769) := X"8FB20024";
		ram_buffer(1770) := X"8FB10020";
		ram_buffer(1771) := X"8FB0001C";
		ram_buffer(1772) := X"03E00008";
		ram_buffer(1773) := X"27BD0040";
		ram_buffer(1774) := X"0C4005AC";
		ram_buffer(1775) := X"02002025";
		ram_buffer(1776) := X"0C400F41";
		ram_buffer(1777) := X"24160001";
		ram_buffer(1778) := X"1000FFD6";
		ram_buffer(1779) := X"00000000";
		ram_buffer(1780) := X"0C4005AC";
		ram_buffer(1781) := X"02002025";
		ram_buffer(1782) := X"0C400F41";
		ram_buffer(1783) := X"00000000";
		ram_buffer(1784) := X"1000FFEA";
		ram_buffer(1785) := X"00001025";
		ram_buffer(1786) := X"3C040100";
		ram_buffer(1787) := X"0C40026D";
		ram_buffer(1788) := X"24845514";
		ram_buffer(1789) := X"1000FF7B";
		ram_buffer(1790) := X"24020002";
		ram_buffer(1791) := X"240502DB";
		ram_buffer(1792) := X"0C40026D";
		ram_buffer(1793) := X"24845514";
		ram_buffer(1794) := X"1000FF7C";
		ram_buffer(1795) := X"00000000";
		ram_buffer(1796) := X"27BDFFE8";
		ram_buffer(1797) := X"00803025";
		ram_buffer(1798) := X"00002825";
		ram_buffer(1799) := X"AFB00010";
		ram_buffer(1800) := X"AFBF0014";
		ram_buffer(1801) := X"0C40061D";
		ram_buffer(1802) := X"24040001";
		ram_buffer(1803) := X"10400009";
		ram_buffer(1804) := X"00408025";
		ram_buffer(1805) := X"AC400004";
		ram_buffer(1806) := X"AC400000";
		ram_buffer(1807) := X"AC40000C";
		ram_buffer(1808) := X"00003825";
		ram_buffer(1809) := X"00003025";
		ram_buffer(1810) := X"00002825";
		ram_buffer(1811) := X"0C40065F";
		ram_buffer(1812) := X"00402025";
		ram_buffer(1813) := X"8FBF0014";
		ram_buffer(1814) := X"02001025";
		ram_buffer(1815) := X"8FB00010";
		ram_buffer(1816) := X"03E00008";
		ram_buffer(1817) := X"27BD0018";
		ram_buffer(1818) := X"27BDFFE0";
		ram_buffer(1819) := X"AFB00010";
		ram_buffer(1820) := X"AFBF001C";
		ram_buffer(1821) := X"AFB20018";
		ram_buffer(1822) := X"AFB10014";
		ram_buffer(1823) := X"14800005";
		ram_buffer(1824) := X"00808025";
		ram_buffer(1825) := X"3C040100";
		ram_buffer(1826) := X"24050241";
		ram_buffer(1827) := X"0C40026D";
		ram_buffer(1828) := X"24845514";
		ram_buffer(1829) := X"8E120004";
		ram_buffer(1830) := X"0C400C4A";
		ram_buffer(1831) := X"00008825";
		ram_buffer(1832) := X"1642000B";
		ram_buffer(1833) := X"00000000";
		ram_buffer(1834) := X"8E02000C";
		ram_buffer(1835) := X"24110001";
		ram_buffer(1836) := X"2442FFFF";
		ram_buffer(1837) := X"14400006";
		ram_buffer(1838) := X"AE02000C";
		ram_buffer(1839) := X"00003825";
		ram_buffer(1840) := X"00003025";
		ram_buffer(1841) := X"00002825";
		ram_buffer(1842) := X"0C40065F";
		ram_buffer(1843) := X"02002025";
		ram_buffer(1844) := X"8FBF001C";
		ram_buffer(1845) := X"02201025";
		ram_buffer(1846) := X"8FB20018";
		ram_buffer(1847) := X"8FB10014";
		ram_buffer(1848) := X"8FB00010";
		ram_buffer(1849) := X"03E00008";
		ram_buffer(1850) := X"27BD0020";
		ram_buffer(1851) := X"27BDFFD0";
		ram_buffer(1852) := X"AFB40024";
		ram_buffer(1853) := X"AFB30020";
		ram_buffer(1854) := X"AFB2001C";
		ram_buffer(1855) := X"AFB00014";
		ram_buffer(1856) := X"AFBF002C";
		ram_buffer(1857) := X"AFB50028";
		ram_buffer(1858) := X"AFB10018";
		ram_buffer(1859) := X"00808025";
		ram_buffer(1860) := X"00A09825";
		ram_buffer(1861) := X"00C0A025";
		ram_buffer(1862) := X"14800005";
		ram_buffer(1863) := X"00E09025";
		ram_buffer(1864) := X"3C040100";
		ram_buffer(1865) := X"2405039F";
		ram_buffer(1866) := X"0C40026D";
		ram_buffer(1867) := X"24845514";
		ram_buffer(1868) := X"16600006";
		ram_buffer(1869) := X"24020002";
		ram_buffer(1870) := X"8E020040";
		ram_buffer(1871) := X"00000000";
		ram_buffer(1872) := X"14400036";
		ram_buffer(1873) := X"240503A0";
		ram_buffer(1874) := X"24020002";
		ram_buffer(1875) := X"16420005";
		ram_buffer(1876) := X"24020001";
		ram_buffer(1877) := X"8E03003C";
		ram_buffer(1878) := X"00000000";
		ram_buffer(1879) := X"14620034";
		ram_buffer(1880) := X"240503A1";
		ram_buffer(1881) := X"8E020038";
		ram_buffer(1882) := X"8E03003C";
		ram_buffer(1883) := X"00000000";
		ram_buffer(1884) := X"0043102B";
		ram_buffer(1885) := X"14400003";
		ram_buffer(1886) := X"24030002";
		ram_buffer(1887) := X"16430018";
		ram_buffer(1888) := X"00000000";
		ram_buffer(1889) := X"92110045";
		ram_buffer(1890) := X"02403025";
		ram_buffer(1891) := X"0011AE00";
		ram_buffer(1892) := X"02602825";
		ram_buffer(1893) := X"0C400556";
		ram_buffer(1894) := X"02002025";
		ram_buffer(1895) := X"0015AE03";
		ram_buffer(1896) := X"2402FFFF";
		ram_buffer(1897) := X"16A20017";
		ram_buffer(1898) := X"00000000";
		ram_buffer(1899) := X"8E020024";
		ram_buffer(1900) := X"00000000";
		ram_buffer(1901) := X"14400003";
		ram_buffer(1902) := X"00000000";
		ram_buffer(1903) := X"10000008";
		ram_buffer(1904) := X"24020001";
		ram_buffer(1905) := X"0C400BB6";
		ram_buffer(1906) := X"26040024";
		ram_buffer(1907) := X"1040FFFB";
		ram_buffer(1908) := X"00000000";
		ram_buffer(1909) := X"12800002";
		ram_buffer(1910) := X"24020001";
		ram_buffer(1911) := X"AE820000";
		ram_buffer(1912) := X"8FBF002C";
		ram_buffer(1913) := X"8FB50028";
		ram_buffer(1914) := X"8FB40024";
		ram_buffer(1915) := X"8FB30020";
		ram_buffer(1916) := X"8FB2001C";
		ram_buffer(1917) := X"8FB10018";
		ram_buffer(1918) := X"8FB00014";
		ram_buffer(1919) := X"03E00008";
		ram_buffer(1920) := X"27BD0030";
		ram_buffer(1921) := X"26310001";
		ram_buffer(1922) := X"00118E00";
		ram_buffer(1923) := X"00118E03";
		ram_buffer(1924) := X"A2110045";
		ram_buffer(1925) := X"1000FFF2";
		ram_buffer(1926) := X"24020001";
		ram_buffer(1927) := X"3C040100";
		ram_buffer(1928) := X"0C40026D";
		ram_buffer(1929) := X"24845514";
		ram_buffer(1930) := X"1000FFC8";
		ram_buffer(1931) := X"24020002";
		ram_buffer(1932) := X"3C040100";
		ram_buffer(1933) := X"0C40026D";
		ram_buffer(1934) := X"24845514";
		ram_buffer(1935) := X"1000FFC9";
		ram_buffer(1936) := X"00000000";
		ram_buffer(1937) := X"27BDFFE0";
		ram_buffer(1938) := X"AFB10018";
		ram_buffer(1939) := X"AFB00014";
		ram_buffer(1940) := X"AFBF001C";
		ram_buffer(1941) := X"00808025";
		ram_buffer(1942) := X"14800005";
		ram_buffer(1943) := X"00A08825";
		ram_buffer(1944) := X"3C040100";
		ram_buffer(1945) := X"2405043C";
		ram_buffer(1946) := X"0C40026D";
		ram_buffer(1947) := X"24845514";
		ram_buffer(1948) := X"8E020040";
		ram_buffer(1949) := X"00000000";
		ram_buffer(1950) := X"10400004";
		ram_buffer(1951) := X"24050440";
		ram_buffer(1952) := X"3C040100";
		ram_buffer(1953) := X"0C40026D";
		ram_buffer(1954) := X"24845514";
		ram_buffer(1955) := X"8E020000";
		ram_buffer(1956) := X"00000000";
		ram_buffer(1957) := X"14400005";
		ram_buffer(1958) := X"00000000";
		ram_buffer(1959) := X"8E020004";
		ram_buffer(1960) := X"00000000";
		ram_buffer(1961) := X"14400026";
		ram_buffer(1962) := X"3C040100";
		ram_buffer(1963) := X"8E030038";
		ram_buffer(1964) := X"8E04003C";
		ram_buffer(1965) := X"00000000";
		ram_buffer(1966) := X"0064202B";
		ram_buffer(1967) := X"10800016";
		ram_buffer(1968) := X"00001025";
		ram_buffer(1969) := X"92020045";
		ram_buffer(1970) := X"24630001";
		ram_buffer(1971) := X"00022600";
		ram_buffer(1972) := X"AE030038";
		ram_buffer(1973) := X"00042603";
		ram_buffer(1974) := X"2403FFFF";
		ram_buffer(1975) := X"14830013";
		ram_buffer(1976) := X"24420001";
		ram_buffer(1977) := X"8E020024";
		ram_buffer(1978) := X"00000000";
		ram_buffer(1979) := X"14400003";
		ram_buffer(1980) := X"00000000";
		ram_buffer(1981) := X"10000008";
		ram_buffer(1982) := X"24020001";
		ram_buffer(1983) := X"0C400BB6";
		ram_buffer(1984) := X"26040024";
		ram_buffer(1985) := X"1040FFFB";
		ram_buffer(1986) := X"00000000";
		ram_buffer(1987) := X"12200002";
		ram_buffer(1988) := X"24020001";
		ram_buffer(1989) := X"AE220000";
		ram_buffer(1990) := X"8FBF001C";
		ram_buffer(1991) := X"8FB10018";
		ram_buffer(1992) := X"8FB00014";
		ram_buffer(1993) := X"03E00008";
		ram_buffer(1994) := X"27BD0020";
		ram_buffer(1995) := X"00021600";
		ram_buffer(1996) := X"00021603";
		ram_buffer(1997) := X"A2020045";
		ram_buffer(1998) := X"1000FFF7";
		ram_buffer(1999) := X"24020001";
		ram_buffer(2000) := X"24050445";
		ram_buffer(2001) := X"0C40026D";
		ram_buffer(2002) := X"24845514";
		ram_buffer(2003) := X"1000FFD7";
		ram_buffer(2004) := X"00000000";
		ram_buffer(2005) := X"27BDFFC8";
		ram_buffer(2006) := X"AFB5002C";
		ram_buffer(2007) := X"AFB30024";
		ram_buffer(2008) := X"AFB00018";
		ram_buffer(2009) := X"AFBF0034";
		ram_buffer(2010) := X"AFB60030";
		ram_buffer(2011) := X"AFB40028";
		ram_buffer(2012) := X"AFB20020";
		ram_buffer(2013) := X"AFB1001C";
		ram_buffer(2014) := X"00808025";
		ram_buffer(2015) := X"00A09825";
		ram_buffer(2016) := X"AFA60040";
		ram_buffer(2017) := X"14800005";
		ram_buffer(2018) := X"00E0A825";
		ram_buffer(2019) := X"3C040100";
		ram_buffer(2020) := X"240504DC";
		ram_buffer(2021) := X"0C40026D";
		ram_buffer(2022) := X"24845514";
		ram_buffer(2023) := X"16600005";
		ram_buffer(2024) := X"00000000";
		ram_buffer(2025) := X"8E020040";
		ram_buffer(2026) := X"00000000";
		ram_buffer(2027) := X"14400096";
		ram_buffer(2028) := X"3C040100";
		ram_buffer(2029) := X"0C400C4D";
		ram_buffer(2030) := X"00000000";
		ram_buffer(2031) := X"14400009";
		ram_buffer(2032) := X"0000B025";
		ram_buffer(2033) := X"8FA20040";
		ram_buffer(2034) := X"00000000";
		ram_buffer(2035) := X"10400005";
		ram_buffer(2036) := X"3C040100";
		ram_buffer(2037) := X"240504E0";
		ram_buffer(2038) := X"0C40026D";
		ram_buffer(2039) := X"24845514";
		ram_buffer(2040) := X"0000B025";
		ram_buffer(2041) := X"2412FFFF";
		ram_buffer(2042) := X"1000004B";
		ram_buffer(2043) := X"26140024";
		ram_buffer(2044) := X"8E020024";
		ram_buffer(2045) := X"AE12000C";
		ram_buffer(2046) := X"10400063";
		ram_buffer(2047) := X"26040024";
		ram_buffer(2048) := X"1000005B";
		ram_buffer(2049) := X"00000000";
		ram_buffer(2050) := X"8FA20040";
		ram_buffer(2051) := X"00000000";
		ram_buffer(2052) := X"14400005";
		ram_buffer(2053) := X"00000000";
		ram_buffer(2054) := X"0C400CE6";
		ram_buffer(2055) := X"00000000";
		ram_buffer(2056) := X"1000005C";
		ram_buffer(2057) := X"00001025";
		ram_buffer(2058) := X"16C00003";
		ram_buffer(2059) := X"00000000";
		ram_buffer(2060) := X"0C400C24";
		ram_buffer(2061) := X"27A40010";
		ram_buffer(2062) := X"0C400CE6";
		ram_buffer(2063) := X"00000000";
		ram_buffer(2064) := X"0C400A98";
		ram_buffer(2065) := X"00000000";
		ram_buffer(2066) := X"0C400CD3";
		ram_buffer(2067) := X"00000000";
		ram_buffer(2068) := X"92020044";
		ram_buffer(2069) := X"00000000";
		ram_buffer(2070) := X"00021600";
		ram_buffer(2071) := X"00021603";
		ram_buffer(2072) := X"14520002";
		ram_buffer(2073) := X"00000000";
		ram_buffer(2074) := X"A2000044";
		ram_buffer(2075) := X"92020045";
		ram_buffer(2076) := X"00000000";
		ram_buffer(2077) := X"00021600";
		ram_buffer(2078) := X"00021603";
		ram_buffer(2079) := X"14520002";
		ram_buffer(2080) := X"00000000";
		ram_buffer(2081) := X"A2000045";
		ram_buffer(2082) := X"0C400CE6";
		ram_buffer(2083) := X"00000000";
		ram_buffer(2084) := X"27A50040";
		ram_buffer(2085) := X"0C4010AC";
		ram_buffer(2086) := X"27A40010";
		ram_buffer(2087) := X"1440004D";
		ram_buffer(2088) := X"00000000";
		ram_buffer(2089) := X"0C400CD3";
		ram_buffer(2090) := X"00000000";
		ram_buffer(2091) := X"8E110038";
		ram_buffer(2092) := X"0C400CE6";
		ram_buffer(2093) := X"00000000";
		ram_buffer(2094) := X"16200040";
		ram_buffer(2095) := X"00000000";
		ram_buffer(2096) := X"8E020000";
		ram_buffer(2097) := X"00000000";
		ram_buffer(2098) := X"14400008";
		ram_buffer(2099) := X"00000000";
		ram_buffer(2100) := X"0C400CD3";
		ram_buffer(2101) := X"00000000";
		ram_buffer(2102) := X"8E040004";
		ram_buffer(2103) := X"0C400C57";
		ram_buffer(2104) := X"00000000";
		ram_buffer(2105) := X"0C400CE6";
		ram_buffer(2106) := X"00000000";
		ram_buffer(2107) := X"8FA50040";
		ram_buffer(2108) := X"0C400B7C";
		ram_buffer(2109) := X"02802025";
		ram_buffer(2110) := X"0C4005AC";
		ram_buffer(2111) := X"02002025";
		ram_buffer(2112) := X"0C400F41";
		ram_buffer(2113) := X"00000000";
		ram_buffer(2114) := X"14400003";
		ram_buffer(2115) := X"24160001";
		ram_buffer(2116) := X"0C400120";
		ram_buffer(2117) := X"00000000";
		ram_buffer(2118) := X"0C400CD3";
		ram_buffer(2119) := X"00000000";
		ram_buffer(2120) := X"8E110038";
		ram_buffer(2121) := X"00000000";
		ram_buffer(2122) := X"1220FFB7";
		ram_buffer(2123) := X"02602825";
		ram_buffer(2124) := X"8E12000C";
		ram_buffer(2125) := X"0C400598";
		ram_buffer(2126) := X"02002025";
		ram_buffer(2127) := X"16A0FFAC";
		ram_buffer(2128) := X"2631FFFF";
		ram_buffer(2129) := X"8E020000";
		ram_buffer(2130) := X"AE110038";
		ram_buffer(2131) := X"14400004";
		ram_buffer(2132) := X"00000000";
		ram_buffer(2133) := X"0C4010F1";
		ram_buffer(2134) := X"00000000";
		ram_buffer(2135) := X"AE020004";
		ram_buffer(2136) := X"8E020010";
		ram_buffer(2137) := X"00000000";
		ram_buffer(2138) := X"10400007";
		ram_buffer(2139) := X"26040010";
		ram_buffer(2140) := X"0C400BB6";
		ram_buffer(2141) := X"00000000";
		ram_buffer(2142) := X"10400003";
		ram_buffer(2143) := X"00000000";
		ram_buffer(2144) := X"0C400120";
		ram_buffer(2145) := X"00000000";
		ram_buffer(2146) := X"0C400CE6";
		ram_buffer(2147) := X"00000000";
		ram_buffer(2148) := X"24020001";
		ram_buffer(2149) := X"8FBF0034";
		ram_buffer(2150) := X"8FB60030";
		ram_buffer(2151) := X"8FB5002C";
		ram_buffer(2152) := X"8FB40028";
		ram_buffer(2153) := X"8FB30024";
		ram_buffer(2154) := X"8FB20020";
		ram_buffer(2155) := X"8FB1001C";
		ram_buffer(2156) := X"8FB00018";
		ram_buffer(2157) := X"03E00008";
		ram_buffer(2158) := X"27BD0038";
		ram_buffer(2159) := X"0C4005AC";
		ram_buffer(2160) := X"02002025";
		ram_buffer(2161) := X"0C400F41";
		ram_buffer(2162) := X"24160001";
		ram_buffer(2163) := X"1000FFD2";
		ram_buffer(2164) := X"00000000";
		ram_buffer(2165) := X"0C4005AC";
		ram_buffer(2166) := X"02002025";
		ram_buffer(2167) := X"0C400F41";
		ram_buffer(2168) := X"00000000";
		ram_buffer(2169) := X"0C400CD3";
		ram_buffer(2170) := X"00000000";
		ram_buffer(2171) := X"8E110038";
		ram_buffer(2172) := X"0C400CE6";
		ram_buffer(2173) := X"00000000";
		ram_buffer(2174) := X"1620FFC7";
		ram_buffer(2175) := X"24160001";
		ram_buffer(2176) := X"1000FFE4";
		ram_buffer(2177) := X"00001025";
		ram_buffer(2178) := X"240504DD";
		ram_buffer(2179) := X"0C40026D";
		ram_buffer(2180) := X"24845514";
		ram_buffer(2181) := X"1000FF67";
		ram_buffer(2182) := X"00000000";
		ram_buffer(2183) := X"27BDFFE0";
		ram_buffer(2184) := X"AFB10014";
		ram_buffer(2185) := X"AFB00010";
		ram_buffer(2186) := X"AFBF001C";
		ram_buffer(2187) := X"AFB20018";
		ram_buffer(2188) := X"00808025";
		ram_buffer(2189) := X"14800005";
		ram_buffer(2190) := X"00A08825";
		ram_buffer(2191) := X"3C040100";
		ram_buffer(2192) := X"24050278";
		ram_buffer(2193) := X"0C40026D";
		ram_buffer(2194) := X"24845514";
		ram_buffer(2195) := X"8E120004";
		ram_buffer(2196) := X"0C400C4A";
		ram_buffer(2197) := X"00000000";
		ram_buffer(2198) := X"1642000C";
		ram_buffer(2199) := X"00003825";
		ram_buffer(2200) := X"8E02000C";
		ram_buffer(2201) := X"00000000";
		ram_buffer(2202) := X"24420001";
		ram_buffer(2203) := X"AE02000C";
		ram_buffer(2204) := X"24020001";
		ram_buffer(2205) := X"8FBF001C";
		ram_buffer(2206) := X"8FB20018";
		ram_buffer(2207) := X"8FB10014";
		ram_buffer(2208) := X"8FB00010";
		ram_buffer(2209) := X"03E00008";
		ram_buffer(2210) := X"27BD0020";
		ram_buffer(2211) := X"02203025";
		ram_buffer(2212) := X"00002825";
		ram_buffer(2213) := X"0C4007D5";
		ram_buffer(2214) := X"02002025";
		ram_buffer(2215) := X"1040FFF5";
		ram_buffer(2216) := X"00000000";
		ram_buffer(2217) := X"8E03000C";
		ram_buffer(2218) := X"00000000";
		ram_buffer(2219) := X"24630001";
		ram_buffer(2220) := X"1000FFF0";
		ram_buffer(2221) := X"AE03000C";
		ram_buffer(2222) := X"27BDFFD0";
		ram_buffer(2223) := X"AFB40024";
		ram_buffer(2224) := X"AFB30020";
		ram_buffer(2225) := X"AFB00014";
		ram_buffer(2226) := X"AFBF002C";
		ram_buffer(2227) := X"AFB50028";
		ram_buffer(2228) := X"AFB2001C";
		ram_buffer(2229) := X"AFB10018";
		ram_buffer(2230) := X"00808025";
		ram_buffer(2231) := X"00A09825";
		ram_buffer(2232) := X"14800005";
		ram_buffer(2233) := X"00C0A025";
		ram_buffer(2234) := X"3C040100";
		ram_buffer(2235) := X"240505A0";
		ram_buffer(2236) := X"0C40026D";
		ram_buffer(2237) := X"24845514";
		ram_buffer(2238) := X"16600005";
		ram_buffer(2239) := X"00000000";
		ram_buffer(2240) := X"8E020040";
		ram_buffer(2241) := X"00000000";
		ram_buffer(2242) := X"1440002C";
		ram_buffer(2243) := X"240505A1";
		ram_buffer(2244) := X"8E120038";
		ram_buffer(2245) := X"00000000";
		ram_buffer(2246) := X"12400019";
		ram_buffer(2247) := X"00001025";
		ram_buffer(2248) := X"92110044";
		ram_buffer(2249) := X"02602825";
		ram_buffer(2250) := X"0011AE00";
		ram_buffer(2251) := X"0C400598";
		ram_buffer(2252) := X"02002025";
		ram_buffer(2253) := X"2652FFFF";
		ram_buffer(2254) := X"0015AE03";
		ram_buffer(2255) := X"2402FFFF";
		ram_buffer(2256) := X"AE120038";
		ram_buffer(2257) := X"16A20017";
		ram_buffer(2258) := X"00000000";
		ram_buffer(2259) := X"8E020010";
		ram_buffer(2260) := X"00000000";
		ram_buffer(2261) := X"14400003";
		ram_buffer(2262) := X"00000000";
		ram_buffer(2263) := X"10000008";
		ram_buffer(2264) := X"24020001";
		ram_buffer(2265) := X"0C400BB6";
		ram_buffer(2266) := X"26040010";
		ram_buffer(2267) := X"1040FFFB";
		ram_buffer(2268) := X"00000000";
		ram_buffer(2269) := X"12800002";
		ram_buffer(2270) := X"24020001";
		ram_buffer(2271) := X"AE820000";
		ram_buffer(2272) := X"8FBF002C";
		ram_buffer(2273) := X"8FB50028";
		ram_buffer(2274) := X"8FB40024";
		ram_buffer(2275) := X"8FB30020";
		ram_buffer(2276) := X"8FB2001C";
		ram_buffer(2277) := X"8FB10018";
		ram_buffer(2278) := X"8FB00014";
		ram_buffer(2279) := X"03E00008";
		ram_buffer(2280) := X"27BD0030";
		ram_buffer(2281) := X"26310001";
		ram_buffer(2282) := X"00118E00";
		ram_buffer(2283) := X"00118E03";
		ram_buffer(2284) := X"A2110044";
		ram_buffer(2285) := X"1000FFF2";
		ram_buffer(2286) := X"24020001";
		ram_buffer(2287) := X"3C040100";
		ram_buffer(2288) := X"0C40026D";
		ram_buffer(2289) := X"24845514";
		ram_buffer(2290) := X"1000FFD1";
		ram_buffer(2291) := X"00000000";
		ram_buffer(2292) := X"27BDFFE0";
		ram_buffer(2293) := X"AFB10014";
		ram_buffer(2294) := X"AFB00010";
		ram_buffer(2295) := X"AFBF001C";
		ram_buffer(2296) := X"AFB20018";
		ram_buffer(2297) := X"00808025";
		ram_buffer(2298) := X"14800005";
		ram_buffer(2299) := X"00A08825";
		ram_buffer(2300) := X"3C040100";
		ram_buffer(2301) := X"240505FC";
		ram_buffer(2302) := X"0C40026D";
		ram_buffer(2303) := X"24845514";
		ram_buffer(2304) := X"16200005";
		ram_buffer(2305) := X"00000000";
		ram_buffer(2306) := X"8E020040";
		ram_buffer(2307) := X"00000000";
		ram_buffer(2308) := X"14400018";
		ram_buffer(2309) := X"240505FD";
		ram_buffer(2310) := X"8E020040";
		ram_buffer(2311) := X"00000000";
		ram_buffer(2312) := X"14400004";
		ram_buffer(2313) := X"240505FE";
		ram_buffer(2314) := X"3C040100";
		ram_buffer(2315) := X"0C40026D";
		ram_buffer(2316) := X"24845514";
		ram_buffer(2317) := X"8E030038";
		ram_buffer(2318) := X"00000000";
		ram_buffer(2319) := X"10600007";
		ram_buffer(2320) := X"00001025";
		ram_buffer(2321) := X"8E12000C";
		ram_buffer(2322) := X"02202825";
		ram_buffer(2323) := X"0C400598";
		ram_buffer(2324) := X"02002025";
		ram_buffer(2325) := X"AE12000C";
		ram_buffer(2326) := X"24020001";
		ram_buffer(2327) := X"8FBF001C";
		ram_buffer(2328) := X"8FB20018";
		ram_buffer(2329) := X"8FB10014";
		ram_buffer(2330) := X"8FB00010";
		ram_buffer(2331) := X"03E00008";
		ram_buffer(2332) := X"27BD0020";
		ram_buffer(2333) := X"3C040100";
		ram_buffer(2334) := X"0C40026D";
		ram_buffer(2335) := X"24845514";
		ram_buffer(2336) := X"1000FFE5";
		ram_buffer(2337) := X"00000000";
		ram_buffer(2338) := X"27BDFFE8";
		ram_buffer(2339) := X"AFB00010";
		ram_buffer(2340) := X"AFBF0014";
		ram_buffer(2341) := X"14800005";
		ram_buffer(2342) := X"00808025";
		ram_buffer(2343) := X"3C040100";
		ram_buffer(2344) := X"2405062F";
		ram_buffer(2345) := X"0C40026D";
		ram_buffer(2346) := X"24845514";
		ram_buffer(2347) := X"0C400CD3";
		ram_buffer(2348) := X"00000000";
		ram_buffer(2349) := X"8E100038";
		ram_buffer(2350) := X"0C400CE6";
		ram_buffer(2351) := X"00000000";
		ram_buffer(2352) := X"8FBF0014";
		ram_buffer(2353) := X"02001025";
		ram_buffer(2354) := X"8FB00010";
		ram_buffer(2355) := X"03E00008";
		ram_buffer(2356) := X"27BD0018";
		ram_buffer(2357) := X"27BDFFE0";
		ram_buffer(2358) := X"AFB10018";
		ram_buffer(2359) := X"AFBF001C";
		ram_buffer(2360) := X"AFB00014";
		ram_buffer(2361) := X"14800005";
		ram_buffer(2362) := X"00808825";
		ram_buffer(2363) := X"3C040100";
		ram_buffer(2364) := X"24050641";
		ram_buffer(2365) := X"0C40026D";
		ram_buffer(2366) := X"24845514";
		ram_buffer(2367) := X"0C400CD3";
		ram_buffer(2368) := X"00000000";
		ram_buffer(2369) := X"8E220038";
		ram_buffer(2370) := X"8E30003C";
		ram_buffer(2371) := X"0C400CE6";
		ram_buffer(2372) := X"02028023";
		ram_buffer(2373) := X"8FBF001C";
		ram_buffer(2374) := X"02001025";
		ram_buffer(2375) := X"8FB10018";
		ram_buffer(2376) := X"8FB00014";
		ram_buffer(2377) := X"03E00008";
		ram_buffer(2378) := X"27BD0020";
		ram_buffer(2379) := X"27BDFFE8";
		ram_buffer(2380) := X"AFB00010";
		ram_buffer(2381) := X"AFBF0014";
		ram_buffer(2382) := X"14800005";
		ram_buffer(2383) := X"00808025";
		ram_buffer(2384) := X"3C040100";
		ram_buffer(2385) := X"24050651";
		ram_buffer(2386) := X"0C40026D";
		ram_buffer(2387) := X"24845514";
		ram_buffer(2388) := X"8FBF0014";
		ram_buffer(2389) := X"8E020038";
		ram_buffer(2390) := X"8FB00010";
		ram_buffer(2391) := X"03E00008";
		ram_buffer(2392) := X"27BD0018";
		ram_buffer(2393) := X"27BDFFE8";
		ram_buffer(2394) := X"AFB00010";
		ram_buffer(2395) := X"AFBF0014";
		ram_buffer(2396) := X"14800005";
		ram_buffer(2397) := X"00808025";
		ram_buffer(2398) := X"3C040100";
		ram_buffer(2399) := X"24050793";
		ram_buffer(2400) := X"0C40026D";
		ram_buffer(2401) := X"24845514";
		ram_buffer(2402) := X"8E020038";
		ram_buffer(2403) := X"8FBF0014";
		ram_buffer(2404) := X"8FB00010";
		ram_buffer(2405) := X"2C420001";
		ram_buffer(2406) := X"03E00008";
		ram_buffer(2407) := X"27BD0018";
		ram_buffer(2408) := X"27BDFFE8";
		ram_buffer(2409) := X"AFB00010";
		ram_buffer(2410) := X"AFBF0014";
		ram_buffer(2411) := X"14800005";
		ram_buffer(2412) := X"00808025";
		ram_buffer(2413) := X"3C040100";
		ram_buffer(2414) := X"240507BA";
		ram_buffer(2415) := X"0C40026D";
		ram_buffer(2416) := X"24845514";
		ram_buffer(2417) := X"8E030038";
		ram_buffer(2418) := X"8E02003C";
		ram_buffer(2419) := X"8FBF0014";
		ram_buffer(2420) := X"00431026";
		ram_buffer(2421) := X"8FB00010";
		ram_buffer(2422) := X"2C420001";
		ram_buffer(2423) := X"03E00008";
		ram_buffer(2424) := X"27BD0018";
		ram_buffer(2425) := X"3C030101";
		ram_buffer(2426) := X"2463596C";
		ram_buffer(2427) := X"00001025";
		ram_buffer(2428) := X"00603025";
		ram_buffer(2429) := X"2407000A";
		ram_buffer(2430) := X"8C680000";
		ram_buffer(2431) := X"00000000";
		ram_buffer(2432) := X"15000007";
		ram_buffer(2433) := X"24420001";
		ram_buffer(2434) := X"2442FFFF";
		ram_buffer(2435) := X"000210C0";
		ram_buffer(2436) := X"00C21021";
		ram_buffer(2437) := X"AC450000";
		ram_buffer(2438) := X"03E00008";
		ram_buffer(2439) := X"AC440004";
		ram_buffer(2440) := X"1447FFF5";
		ram_buffer(2441) := X"24630008";
		ram_buffer(2442) := X"03E00008";
		ram_buffer(2443) := X"00000000";
		ram_buffer(2444) := X"3C030101";
		ram_buffer(2445) := X"2463596C";
		ram_buffer(2446) := X"00001025";
		ram_buffer(2447) := X"00602825";
		ram_buffer(2448) := X"2406000A";
		ram_buffer(2449) := X"8C670004";
		ram_buffer(2450) := X"00000000";
		ram_buffer(2451) := X"14E40007";
		ram_buffer(2452) := X"24420001";
		ram_buffer(2453) := X"2442FFFF";
		ram_buffer(2454) := X"000210C0";
		ram_buffer(2455) := X"00A21021";
		ram_buffer(2456) := X"8C420000";
		ram_buffer(2457) := X"03E00008";
		ram_buffer(2458) := X"00000000";
		ram_buffer(2459) := X"1446FFF5";
		ram_buffer(2460) := X"24630008";
		ram_buffer(2461) := X"03E00008";
		ram_buffer(2462) := X"00001025";
		ram_buffer(2463) := X"3C030101";
		ram_buffer(2464) := X"2463596C";
		ram_buffer(2465) := X"00001025";
		ram_buffer(2466) := X"00602825";
		ram_buffer(2467) := X"2406000A";
		ram_buffer(2468) := X"8C670004";
		ram_buffer(2469) := X"00000000";
		ram_buffer(2470) := X"14E40007";
		ram_buffer(2471) := X"24420001";
		ram_buffer(2472) := X"2442FFFF";
		ram_buffer(2473) := X"000210C0";
		ram_buffer(2474) := X"00A21021";
		ram_buffer(2475) := X"AC400000";
		ram_buffer(2476) := X"03E00008";
		ram_buffer(2477) := X"AC400004";
		ram_buffer(2478) := X"1446FFF5";
		ram_buffer(2479) := X"24630008";
		ram_buffer(2480) := X"03E00008";
		ram_buffer(2481) := X"00000000";
		ram_buffer(2482) := X"27BDFFE8";
		ram_buffer(2483) := X"AFB00010";
		ram_buffer(2484) := X"AFBF0014";
		ram_buffer(2485) := X"14800005";
		ram_buffer(2486) := X"00808025";
		ram_buffer(2487) := X"3C040100";
		ram_buffer(2488) := X"2405065D";
		ram_buffer(2489) := X"0C40026D";
		ram_buffer(2490) := X"24845514";
		ram_buffer(2491) := X"0C40099F";
		ram_buffer(2492) := X"02002025";
		ram_buffer(2493) := X"8FBF0014";
		ram_buffer(2494) := X"02002025";
		ram_buffer(2495) := X"8FB00010";
		ram_buffer(2496) := X"0840135A";
		ram_buffer(2497) := X"27BD0018";
		ram_buffer(2498) := X"8C820000";
		ram_buffer(2499) := X"00000000";
		ram_buffer(2500) := X"10400027";
		ram_buffer(2501) := X"24870008";
		ram_buffer(2502) := X"8C820004";
		ram_buffer(2503) := X"00000000";
		ram_buffer(2504) := X"8C420004";
		ram_buffer(2505) := X"00000000";
		ram_buffer(2506) := X"14470004";
		ram_buffer(2507) := X"AC820004";
		ram_buffer(2508) := X"8C82000C";
		ram_buffer(2509) := X"00000000";
		ram_buffer(2510) := X"AC820004";
		ram_buffer(2511) := X"8C820004";
		ram_buffer(2512) := X"00000000";
		ram_buffer(2513) := X"8C49000C";
		ram_buffer(2514) := X"8C820004";
		ram_buffer(2515) := X"00000000";
		ram_buffer(2516) := X"8C420004";
		ram_buffer(2517) := X"00000000";
		ram_buffer(2518) := X"14E20004";
		ram_buffer(2519) := X"AC820004";
		ram_buffer(2520) := X"8C82000C";
		ram_buffer(2521) := X"00000000";
		ram_buffer(2522) := X"AC820004";
		ram_buffer(2523) := X"8C820004";
		ram_buffer(2524) := X"00A03025";
		ram_buffer(2525) := X"8C42000C";
		ram_buffer(2526) := X"00000000";
		ram_buffer(2527) := X"24430034";
		ram_buffer(2528) := X"244A0044";
		ram_buffer(2529) := X"806B0000";
		ram_buffer(2530) := X"80C80000";
		ram_buffer(2531) := X"00000000";
		ram_buffer(2532) := X"150B0005";
		ram_buffer(2533) := X"00000000";
		ram_buffer(2534) := X"11000006";
		ram_buffer(2535) := X"24630001";
		ram_buffer(2536) := X"146AFFF8";
		ram_buffer(2537) := X"24C60001";
		ram_buffer(2538) := X"1522FFE7";
		ram_buffer(2539) := X"00000000";
		ram_buffer(2540) := X"00001025";
		ram_buffer(2541) := X"03E00008";
		ram_buffer(2542) := X"00000000";
		ram_buffer(2543) := X"8F828050";
		ram_buffer(2544) := X"00000000";
		ram_buffer(2545) := X"8C420000";
		ram_buffer(2546) := X"00000000";
		ram_buffer(2547) := X"14400005";
		ram_buffer(2548) := X"00000000";
		ram_buffer(2549) := X"2402FFFF";
		ram_buffer(2550) := X"AF828024";
		ram_buffer(2551) := X"03E00008";
		ram_buffer(2552) := X"00000000";
		ram_buffer(2553) := X"8F828050";
		ram_buffer(2554) := X"00000000";
		ram_buffer(2555) := X"8C42000C";
		ram_buffer(2556) := X"00000000";
		ram_buffer(2557) := X"8C42000C";
		ram_buffer(2558) := X"00000000";
		ram_buffer(2559) := X"8C420004";
		ram_buffer(2560) := X"1000FFF5";
		ram_buffer(2561) := X"00000000";
		ram_buffer(2562) := X"27BDFFE8";
		ram_buffer(2563) := X"AFB00010";
		ram_buffer(2564) := X"AFBF0014";
		ram_buffer(2565) := X"14800005";
		ram_buffer(2566) := X"00808025";
		ram_buffer(2567) := X"3C040100";
		ram_buffer(2568) := X"24050688";
		ram_buffer(2569) := X"0C40026D";
		ram_buffer(2570) := X"2484552C";
		ram_buffer(2571) := X"3C030100";
		ram_buffer(2572) := X"8E040014";
		ram_buffer(2573) := X"24635630";
		ram_buffer(2574) := X"14830007";
		ram_buffer(2575) := X"00001025";
		ram_buffer(2576) := X"3C030100";
		ram_buffer(2577) := X"8E040028";
		ram_buffer(2578) := X"24635658";
		ram_buffer(2579) := X"10830002";
		ram_buffer(2580) := X"00000000";
		ram_buffer(2581) := X"2C820001";
		ram_buffer(2582) := X"8FBF0014";
		ram_buffer(2583) := X"8FB00010";
		ram_buffer(2584) := X"03E00008";
		ram_buffer(2585) := X"27BD0018";
		ram_buffer(2586) := X"27BDFFE0";
		ram_buffer(2587) := X"AFB10014";
		ram_buffer(2588) := X"AFB00010";
		ram_buffer(2589) := X"8F918040";
		ram_buffer(2590) := X"00808025";
		ram_buffer(2591) := X"8F828018";
		ram_buffer(2592) := X"8F848018";
		ram_buffer(2593) := X"AFB20018";
		ram_buffer(2594) := X"AFBF001C";
		ram_buffer(2595) := X"24840004";
		ram_buffer(2596) := X"A0400055";
		ram_buffer(2597) := X"0C400545";
		ram_buffer(2598) := X"00A09025";
		ram_buffer(2599) := X"2402FFFF";
		ram_buffer(2600) := X"1602000D";
		ram_buffer(2601) := X"00000000";
		ram_buffer(2602) := X"1240000C";
		ram_buffer(2603) := X"02308021";
		ram_buffer(2604) := X"8F858018";
		ram_buffer(2605) := X"8FBF001C";
		ram_buffer(2606) := X"8FB20018";
		ram_buffer(2607) := X"8FB10014";
		ram_buffer(2608) := X"8FB00010";
		ram_buffer(2609) := X"3C040100";
		ram_buffer(2610) := X"24A50004";
		ram_buffer(2611) := X"24845630";
		ram_buffer(2612) := X"0840051C";
		ram_buffer(2613) := X"27BD0020";
		ram_buffer(2614) := X"02308021";
		ram_buffer(2615) := X"8F828018";
		ram_buffer(2616) := X"0211882B";
		ram_buffer(2617) := X"1220000A";
		ram_buffer(2618) := X"AC500004";
		ram_buffer(2619) := X"8F84804C";
		ram_buffer(2620) := X"8F858018";
		ram_buffer(2621) := X"8FBF001C";
		ram_buffer(2622) := X"8FB20018";
		ram_buffer(2623) := X"8FB10014";
		ram_buffer(2624) := X"8FB00010";
		ram_buffer(2625) := X"24A50004";
		ram_buffer(2626) := X"0840052A";
		ram_buffer(2627) := X"27BD0020";
		ram_buffer(2628) := X"8F848050";
		ram_buffer(2629) := X"8F858018";
		ram_buffer(2630) := X"0C40052A";
		ram_buffer(2631) := X"24A50004";
		ram_buffer(2632) := X"8F828024";
		ram_buffer(2633) := X"00000000";
		ram_buffer(2634) := X"0202102B";
		ram_buffer(2635) := X"10400002";
		ram_buffer(2636) := X"00000000";
		ram_buffer(2637) := X"AF908024";
		ram_buffer(2638) := X"8FBF001C";
		ram_buffer(2639) := X"8FB20018";
		ram_buffer(2640) := X"8FB10014";
		ram_buffer(2641) := X"8FB00010";
		ram_buffer(2642) := X"03E00008";
		ram_buffer(2643) := X"27BD0020";
		ram_buffer(2644) := X"14800003";
		ram_buffer(2645) := X"00000000";
		ram_buffer(2646) := X"8F848018";
		ram_buffer(2647) := X"00000000";
		ram_buffer(2648) := X"8C82002C";
		ram_buffer(2649) := X"03E00008";
		ram_buffer(2650) := X"00000000";
		ram_buffer(2651) := X"27BDFFE0";
		ram_buffer(2652) := X"AFB10014";
		ram_buffer(2653) := X"AFBF001C";
		ram_buffer(2654) := X"AFB20018";
		ram_buffer(2655) := X"AFB00010";
		ram_buffer(2656) := X"14800005";
		ram_buffer(2657) := X"00808825";
		ram_buffer(2658) := X"3C040100";
		ram_buffer(2659) := X"240506E9";
		ram_buffer(2660) := X"0C40026D";
		ram_buffer(2661) := X"2484552C";
		ram_buffer(2662) := X"0C400A02";
		ram_buffer(2663) := X"02202025";
		ram_buffer(2664) := X"1040001C";
		ram_buffer(2665) := X"00008025";
		ram_buffer(2666) := X"8F82801C";
		ram_buffer(2667) := X"00000000";
		ram_buffer(2668) := X"1440001F";
		ram_buffer(2669) := X"3C040100";
		ram_buffer(2670) := X"8F828018";
		ram_buffer(2671) := X"8E30002C";
		ram_buffer(2672) := X"8C42002C";
		ram_buffer(2673) := X"26320004";
		ram_buffer(2674) := X"02402025";
		ram_buffer(2675) := X"0C400545";
		ram_buffer(2676) := X"0202802B";
		ram_buffer(2677) := X"8E24002C";
		ram_buffer(2678) := X"8F82803C";
		ram_buffer(2679) := X"00000000";
		ram_buffer(2680) := X"0044102B";
		ram_buffer(2681) := X"10400002";
		ram_buffer(2682) := X"3A100001";
		ram_buffer(2683) := X"AF84803C";
		ram_buffer(2684) := X"00041080";
		ram_buffer(2685) := X"00441021";
		ram_buffer(2686) := X"3C040100";
		ram_buffer(2687) := X"00021080";
		ram_buffer(2688) := X"24845694";
		ram_buffer(2689) := X"02402825";
		ram_buffer(2690) := X"00822021";
		ram_buffer(2691) := X"0C40051C";
		ram_buffer(2692) := X"00000000";
		ram_buffer(2693) := X"8FBF001C";
		ram_buffer(2694) := X"02001025";
		ram_buffer(2695) := X"8FB20018";
		ram_buffer(2696) := X"8FB10014";
		ram_buffer(2697) := X"8FB00010";
		ram_buffer(2698) := X"03E00008";
		ram_buffer(2699) := X"27BD0020";
		ram_buffer(2700) := X"26250018";
		ram_buffer(2701) := X"1000FFF5";
		ram_buffer(2702) := X"24845658";
		ram_buffer(2703) := X"27BDFFE8";
		ram_buffer(2704) := X"AFBF0014";
		ram_buffer(2705) := X"0C400284";
		ram_buffer(2706) := X"00000000";
		ram_buffer(2707) := X"8FBF0014";
		ram_buffer(2708) := X"27BD0018";
		ram_buffer(2709) := X"AF808038";
		ram_buffer(2710) := X"084012C0";
		ram_buffer(2711) := X"00000000";
		ram_buffer(2712) := X"8F82801C";
		ram_buffer(2713) := X"00000000";
		ram_buffer(2714) := X"24420001";
		ram_buffer(2715) := X"AF82801C";
		ram_buffer(2716) := X"03E00008";
		ram_buffer(2717) := X"00000000";
		ram_buffer(2718) := X"8F828040";
		ram_buffer(2719) := X"03E00008";
		ram_buffer(2720) := X"00000000";
		ram_buffer(2721) := X"8F828040";
		ram_buffer(2722) := X"03E00008";
		ram_buffer(2723) := X"00000000";
		ram_buffer(2724) := X"8F828044";
		ram_buffer(2725) := X"03E00008";
		ram_buffer(2726) := X"00000000";
		ram_buffer(2727) := X"27BDFFE8";
		ram_buffer(2728) := X"AFB00010";
		ram_buffer(2729) := X"AFBF0014";
		ram_buffer(2730) := X"14800008";
		ram_buffer(2731) := X"00808025";
		ram_buffer(2732) := X"8F908018";
		ram_buffer(2733) := X"00000000";
		ram_buffer(2734) := X"16000004";
		ram_buffer(2735) := X"24050893";
		ram_buffer(2736) := X"3C040100";
		ram_buffer(2737) := X"0C40026D";
		ram_buffer(2738) := X"2484552C";
		ram_buffer(2739) := X"8FBF0014";
		ram_buffer(2740) := X"26020034";
		ram_buffer(2741) := X"8FB00010";
		ram_buffer(2742) := X"03E00008";
		ram_buffer(2743) := X"27BD0018";
		ram_buffer(2744) := X"8F828020";
		ram_buffer(2745) := X"27BDFFE8";
		ram_buffer(2746) := X"14400005";
		ram_buffer(2747) := X"AFBF0014";
		ram_buffer(2748) := X"3C040100";
		ram_buffer(2749) := X"24050966";
		ram_buffer(2750) := X"0C40026D";
		ram_buffer(2751) := X"2484552C";
		ram_buffer(2752) := X"8FBF0014";
		ram_buffer(2753) := X"8F828020";
		ram_buffer(2754) := X"03E00008";
		ram_buffer(2755) := X"27BD0018";
		ram_buffer(2756) := X"8F82801C";
		ram_buffer(2757) := X"27BDFFD8";
		ram_buffer(2758) := X"AFBF0024";
		ram_buffer(2759) := X"AFB40020";
		ram_buffer(2760) := X"AFB3001C";
		ram_buffer(2761) := X"AFB20018";
		ram_buffer(2762) := X"AFB10014";
		ram_buffer(2763) := X"1440006D";
		ram_buffer(2764) := X"AFB00010";
		ram_buffer(2765) := X"8F918040";
		ram_buffer(2766) := X"00000000";
		ram_buffer(2767) := X"26310001";
		ram_buffer(2768) := X"AF918040";
		ram_buffer(2769) := X"16200015";
		ram_buffer(2770) := X"00000000";
		ram_buffer(2771) := X"8F828050";
		ram_buffer(2772) := X"00000000";
		ram_buffer(2773) := X"8C420000";
		ram_buffer(2774) := X"00000000";
		ram_buffer(2775) := X"10400004";
		ram_buffer(2776) := X"240509E4";
		ram_buffer(2777) := X"3C040100";
		ram_buffer(2778) := X"0C40026D";
		ram_buffer(2779) := X"2484552C";
		ram_buffer(2780) := X"8F828050";
		ram_buffer(2781) := X"8F83804C";
		ram_buffer(2782) := X"00000000";
		ram_buffer(2783) := X"AF838050";
		ram_buffer(2784) := X"AF82804C";
		ram_buffer(2785) := X"8F82802C";
		ram_buffer(2786) := X"00000000";
		ram_buffer(2787) := X"24420001";
		ram_buffer(2788) := X"AF82802C";
		ram_buffer(2789) := X"0C4009EF";
		ram_buffer(2790) := X"00000000";
		ram_buffer(2791) := X"8F828024";
		ram_buffer(2792) := X"3C100100";
		ram_buffer(2793) := X"0222102B";
		ram_buffer(2794) := X"26105694";
		ram_buffer(2795) := X"14400008";
		ram_buffer(2796) := X"00009825";
		ram_buffer(2797) := X"8F828050";
		ram_buffer(2798) := X"00000000";
		ram_buffer(2799) := X"8C420000";
		ram_buffer(2800) := X"00000000";
		ram_buffer(2801) := X"1440001E";
		ram_buffer(2802) := X"2402FFFF";
		ram_buffer(2803) := X"AF828024";
		ram_buffer(2804) := X"8F828018";
		ram_buffer(2805) := X"00000000";
		ram_buffer(2806) := X"8C43002C";
		ram_buffer(2807) := X"00000000";
		ram_buffer(2808) := X"00031080";
		ram_buffer(2809) := X"00431021";
		ram_buffer(2810) := X"00021080";
		ram_buffer(2811) := X"02028021";
		ram_buffer(2812) := X"8E020000";
		ram_buffer(2813) := X"00000000";
		ram_buffer(2814) := X"2C420002";
		ram_buffer(2815) := X"14400002";
		ram_buffer(2816) := X"00000000";
		ram_buffer(2817) := X"24130001";
		ram_buffer(2818) := X"8F828030";
		ram_buffer(2819) := X"00000000";
		ram_buffer(2820) := X"10400002";
		ram_buffer(2821) := X"00000000";
		ram_buffer(2822) := X"24130001";
		ram_buffer(2823) := X"8FBF0024";
		ram_buffer(2824) := X"02601025";
		ram_buffer(2825) := X"8FB40020";
		ram_buffer(2826) := X"8FB3001C";
		ram_buffer(2827) := X"8FB20018";
		ram_buffer(2828) := X"8FB10014";
		ram_buffer(2829) := X"8FB00010";
		ram_buffer(2830) := X"03E00008";
		ram_buffer(2831) := X"27BD0028";
		ram_buffer(2832) := X"8F828050";
		ram_buffer(2833) := X"00000000";
		ram_buffer(2834) := X"8C42000C";
		ram_buffer(2835) := X"00000000";
		ram_buffer(2836) := X"8C52000C";
		ram_buffer(2837) := X"00000000";
		ram_buffer(2838) := X"8E420004";
		ram_buffer(2839) := X"00000000";
		ram_buffer(2840) := X"0222182B";
		ram_buffer(2841) := X"1460FFD9";
		ram_buffer(2842) := X"26540004";
		ram_buffer(2843) := X"0C400545";
		ram_buffer(2844) := X"02802025";
		ram_buffer(2845) := X"8E420028";
		ram_buffer(2846) := X"00000000";
		ram_buffer(2847) := X"10400003";
		ram_buffer(2848) := X"00000000";
		ram_buffer(2849) := X"0C400545";
		ram_buffer(2850) := X"26440018";
		ram_buffer(2851) := X"8E42002C";
		ram_buffer(2852) := X"8F83803C";
		ram_buffer(2853) := X"00000000";
		ram_buffer(2854) := X"0062182B";
		ram_buffer(2855) := X"10600002";
		ram_buffer(2856) := X"00000000";
		ram_buffer(2857) := X"AF82803C";
		ram_buffer(2858) := X"00022080";
		ram_buffer(2859) := X"00822021";
		ram_buffer(2860) := X"00042080";
		ram_buffer(2861) := X"02802825";
		ram_buffer(2862) := X"0C40051C";
		ram_buffer(2863) := X"02042021";
		ram_buffer(2864) := X"8F838018";
		ram_buffer(2865) := X"8E42002C";
		ram_buffer(2866) := X"8C63002C";
		ram_buffer(2867) := X"00000000";
		ram_buffer(2868) := X"0043102B";
		ram_buffer(2869) := X"1440FFB7";
		ram_buffer(2870) := X"00000000";
		ram_buffer(2871) := X"1000FFB5";
		ram_buffer(2872) := X"24130001";
		ram_buffer(2873) := X"8F828034";
		ram_buffer(2874) := X"00009825";
		ram_buffer(2875) := X"24420001";
		ram_buffer(2876) := X"AF828034";
		ram_buffer(2877) := X"1000FFC4";
		ram_buffer(2878) := X"00000000";
		ram_buffer(2879) := X"8F82801C";
		ram_buffer(2880) := X"27BDFFD8";
		ram_buffer(2881) := X"AFBF0024";
		ram_buffer(2882) := X"AFB30020";
		ram_buffer(2883) := X"AFB2001C";
		ram_buffer(2884) := X"AFB10018";
		ram_buffer(2885) := X"1040000A";
		ram_buffer(2886) := X"AFB00014";
		ram_buffer(2887) := X"24020001";
		ram_buffer(2888) := X"AF828030";
		ram_buffer(2889) := X"8FBF0024";
		ram_buffer(2890) := X"8FB30020";
		ram_buffer(2891) := X"8FB2001C";
		ram_buffer(2892) := X"8FB10018";
		ram_buffer(2893) := X"8FB00014";
		ram_buffer(2894) := X"03E00008";
		ram_buffer(2895) := X"27BD0028";
		ram_buffer(2896) := X"AF808030";
		ram_buffer(2897) := X"8F90803C";
		ram_buffer(2898) := X"3C120100";
		ram_buffer(2899) := X"00108880";
		ram_buffer(2900) := X"02308821";
		ram_buffer(2901) := X"00118880";
		ram_buffer(2902) := X"26525694";
		ram_buffer(2903) := X"3C130100";
		ram_buffer(2904) := X"02518821";
		ram_buffer(2905) := X"2673552C";
		ram_buffer(2906) := X"8E220000";
		ram_buffer(2907) := X"00000000";
		ram_buffer(2908) := X"10400018";
		ram_buffer(2909) := X"00101880";
		ram_buffer(2910) := X"00701021";
		ram_buffer(2911) := X"00021080";
		ram_buffer(2912) := X"02422021";
		ram_buffer(2913) := X"8C850004";
		ram_buffer(2914) := X"24420008";
		ram_buffer(2915) := X"8CA50004";
		ram_buffer(2916) := X"02421021";
		ram_buffer(2917) := X"14A20004";
		ram_buffer(2918) := X"AC850004";
		ram_buffer(2919) := X"8CA20004";
		ram_buffer(2920) := X"00000000";
		ram_buffer(2921) := X"AC820004";
		ram_buffer(2922) := X"00701821";
		ram_buffer(2923) := X"00031880";
		ram_buffer(2924) := X"02439021";
		ram_buffer(2925) := X"8E420004";
		ram_buffer(2926) := X"00000000";
		ram_buffer(2927) := X"8C42000C";
		ram_buffer(2928) := X"00000000";
		ram_buffer(2929) := X"AF828018";
		ram_buffer(2930) := X"AF90803C";
		ram_buffer(2931) := X"1000FFD5";
		ram_buffer(2932) := X"00000000";
		ram_buffer(2933) := X"16000003";
		ram_buffer(2934) := X"24050B05";
		ram_buffer(2935) := X"0C40026D";
		ram_buffer(2936) := X"02602025";
		ram_buffer(2937) := X"2610FFFF";
		ram_buffer(2938) := X"1000FFDF";
		ram_buffer(2939) := X"2631FFEC";
		ram_buffer(2940) := X"27BDFFE0";
		ram_buffer(2941) := X"AFB10018";
		ram_buffer(2942) := X"AFB00014";
		ram_buffer(2943) := X"AFBF001C";
		ram_buffer(2944) := X"00808025";
		ram_buffer(2945) := X"14800005";
		ram_buffer(2946) := X"00A08825";
		ram_buffer(2947) := X"3C040100";
		ram_buffer(2948) := X"24050B15";
		ram_buffer(2949) := X"0C40026D";
		ram_buffer(2950) := X"2484552C";
		ram_buffer(2951) := X"8F858018";
		ram_buffer(2952) := X"02002025";
		ram_buffer(2953) := X"0C40052A";
		ram_buffer(2954) := X"24A50018";
		ram_buffer(2955) := X"8FBF001C";
		ram_buffer(2956) := X"8FB00014";
		ram_buffer(2957) := X"02202025";
		ram_buffer(2958) := X"8FB10018";
		ram_buffer(2959) := X"24050001";
		ram_buffer(2960) := X"08400A1A";
		ram_buffer(2961) := X"27BD0020";
		ram_buffer(2962) := X"27BDFFE0";
		ram_buffer(2963) := X"AFB20018";
		ram_buffer(2964) := X"AFB10014";
		ram_buffer(2965) := X"AFB00010";
		ram_buffer(2966) := X"AFBF001C";
		ram_buffer(2967) := X"00808825";
		ram_buffer(2968) := X"00A08025";
		ram_buffer(2969) := X"14800005";
		ram_buffer(2970) := X"00C09025";
		ram_buffer(2971) := X"3C040100";
		ram_buffer(2972) := X"24050B26";
		ram_buffer(2973) := X"0C40026D";
		ram_buffer(2974) := X"2484552C";
		ram_buffer(2975) := X"8F82801C";
		ram_buffer(2976) := X"00000000";
		ram_buffer(2977) := X"14400004";
		ram_buffer(2978) := X"3C040100";
		ram_buffer(2979) := X"24050B2A";
		ram_buffer(2980) := X"0C40026D";
		ram_buffer(2981) := X"2484552C";
		ram_buffer(2982) := X"8F828018";
		ram_buffer(2983) := X"3C038000";
		ram_buffer(2984) := X"8F858018";
		ram_buffer(2985) := X"02038025";
		ram_buffer(2986) := X"02202025";
		ram_buffer(2987) := X"AC500018";
		ram_buffer(2988) := X"0C40051C";
		ram_buffer(2989) := X"24A50018";
		ram_buffer(2990) := X"8FBF001C";
		ram_buffer(2991) := X"8FB10014";
		ram_buffer(2992) := X"8FB00010";
		ram_buffer(2993) := X"02402025";
		ram_buffer(2994) := X"8FB20018";
		ram_buffer(2995) := X"24050001";
		ram_buffer(2996) := X"08400A1A";
		ram_buffer(2997) := X"27BD0020";
		ram_buffer(2998) := X"8C82000C";
		ram_buffer(2999) := X"27BDFFE0";
		ram_buffer(3000) := X"AFB00014";
		ram_buffer(3001) := X"8C50000C";
		ram_buffer(3002) := X"AFBF001C";
		ram_buffer(3003) := X"16000005";
		ram_buffer(3004) := X"AFB10018";
		ram_buffer(3005) := X"3C040100";
		ram_buffer(3006) := X"24050B70";
		ram_buffer(3007) := X"0C40026D";
		ram_buffer(3008) := X"2484552C";
		ram_buffer(3009) := X"26110018";
		ram_buffer(3010) := X"0C400545";
		ram_buffer(3011) := X"02202025";
		ram_buffer(3012) := X"8F82801C";
		ram_buffer(3013) := X"00000000";
		ram_buffer(3014) := X"14400022";
		ram_buffer(3015) := X"3C040100";
		ram_buffer(3016) := X"26110004";
		ram_buffer(3017) := X"0C400545";
		ram_buffer(3018) := X"02202025";
		ram_buffer(3019) := X"8E04002C";
		ram_buffer(3020) := X"8F82803C";
		ram_buffer(3021) := X"00000000";
		ram_buffer(3022) := X"0044102B";
		ram_buffer(3023) := X"10400002";
		ram_buffer(3024) := X"00000000";
		ram_buffer(3025) := X"AF84803C";
		ram_buffer(3026) := X"00041080";
		ram_buffer(3027) := X"00441021";
		ram_buffer(3028) := X"3C040100";
		ram_buffer(3029) := X"00021080";
		ram_buffer(3030) := X"24845694";
		ram_buffer(3031) := X"02202825";
		ram_buffer(3032) := X"00822021";
		ram_buffer(3033) := X"0C40051C";
		ram_buffer(3034) := X"00000000";
		ram_buffer(3035) := X"8F828018";
		ram_buffer(3036) := X"8E03002C";
		ram_buffer(3037) := X"8C42002C";
		ram_buffer(3038) := X"00000000";
		ram_buffer(3039) := X"0043182B";
		ram_buffer(3040) := X"10600003";
		ram_buffer(3041) := X"00001025";
		ram_buffer(3042) := X"24020001";
		ram_buffer(3043) := X"AF828030";
		ram_buffer(3044) := X"8FBF001C";
		ram_buffer(3045) := X"8FB10018";
		ram_buffer(3046) := X"8FB00014";
		ram_buffer(3047) := X"03E00008";
		ram_buffer(3048) := X"27BD0020";
		ram_buffer(3049) := X"02202825";
		ram_buffer(3050) := X"1000FFEE";
		ram_buffer(3051) := X"24845658";
		ram_buffer(3052) := X"8F82801C";
		ram_buffer(3053) := X"27BDFFE0";
		ram_buffer(3054) := X"AFB10018";
		ram_buffer(3055) := X"AFB00014";
		ram_buffer(3056) := X"AFBF001C";
		ram_buffer(3057) := X"00808825";
		ram_buffer(3058) := X"14400005";
		ram_buffer(3059) := X"00A08025";
		ram_buffer(3060) := X"3C040100";
		ram_buffer(3061) := X"24050BA8";
		ram_buffer(3062) := X"0C40026D";
		ram_buffer(3063) := X"2484552C";
		ram_buffer(3064) := X"3C028000";
		ram_buffer(3065) := X"02028025";
		ram_buffer(3066) := X"AE300000";
		ram_buffer(3067) := X"8E30000C";
		ram_buffer(3068) := X"00000000";
		ram_buffer(3069) := X"16000004";
		ram_buffer(3070) := X"24050BB0";
		ram_buffer(3071) := X"3C040100";
		ram_buffer(3072) := X"0C40026D";
		ram_buffer(3073) := X"2484552C";
		ram_buffer(3074) := X"02202025";
		ram_buffer(3075) := X"0C400545";
		ram_buffer(3076) := X"26110004";
		ram_buffer(3077) := X"0C400545";
		ram_buffer(3078) := X"02202025";
		ram_buffer(3079) := X"8E04002C";
		ram_buffer(3080) := X"8F82803C";
		ram_buffer(3081) := X"00000000";
		ram_buffer(3082) := X"0044102B";
		ram_buffer(3083) := X"10400002";
		ram_buffer(3084) := X"00000000";
		ram_buffer(3085) := X"AF84803C";
		ram_buffer(3086) := X"00041080";
		ram_buffer(3087) := X"00441021";
		ram_buffer(3088) := X"3C040100";
		ram_buffer(3089) := X"00021080";
		ram_buffer(3090) := X"24845694";
		ram_buffer(3091) := X"00822021";
		ram_buffer(3092) := X"0C40051C";
		ram_buffer(3093) := X"02202825";
		ram_buffer(3094) := X"8F828018";
		ram_buffer(3095) := X"8E03002C";
		ram_buffer(3096) := X"8C42002C";
		ram_buffer(3097) := X"00000000";
		ram_buffer(3098) := X"0043182B";
		ram_buffer(3099) := X"10600003";
		ram_buffer(3100) := X"00001025";
		ram_buffer(3101) := X"24020001";
		ram_buffer(3102) := X"AF828030";
		ram_buffer(3103) := X"8FBF001C";
		ram_buffer(3104) := X"8FB10018";
		ram_buffer(3105) := X"8FB00014";
		ram_buffer(3106) := X"03E00008";
		ram_buffer(3107) := X"27BD0020";
		ram_buffer(3108) := X"27BDFFE8";
		ram_buffer(3109) := X"AFB00010";
		ram_buffer(3110) := X"AFBF0014";
		ram_buffer(3111) := X"14800005";
		ram_buffer(3112) := X"00808025";
		ram_buffer(3113) := X"3C040100";
		ram_buffer(3114) := X"24050BD0";
		ram_buffer(3115) := X"0C40026D";
		ram_buffer(3116) := X"2484552C";
		ram_buffer(3117) := X"8F82802C";
		ram_buffer(3118) := X"8FBF0014";
		ram_buffer(3119) := X"AE020000";
		ram_buffer(3120) := X"8F828040";
		ram_buffer(3121) := X"00000000";
		ram_buffer(3122) := X"AE020004";
		ram_buffer(3123) := X"8FB00010";
		ram_buffer(3124) := X"03E00008";
		ram_buffer(3125) := X"27BD0018";
		ram_buffer(3126) := X"24020001";
		ram_buffer(3127) := X"AF828030";
		ram_buffer(3128) := X"03E00008";
		ram_buffer(3129) := X"00000000";
		ram_buffer(3130) := X"14800003";
		ram_buffer(3131) := X"00000000";
		ram_buffer(3132) := X"8F848018";
		ram_buffer(3133) := X"00000000";
		ram_buffer(3134) := X"8C840030";
		ram_buffer(3135) := X"240500A5";
		ram_buffer(3136) := X"00801825";
		ram_buffer(3137) := X"90660000";
		ram_buffer(3138) := X"00000000";
		ram_buffer(3139) := X"10C50004";
		ram_buffer(3140) := X"00641023";
		ram_buffer(3141) := X"00021082";
		ram_buffer(3142) := X"03E00008";
		ram_buffer(3143) := X"3042FFFF";
		ram_buffer(3144) := X"1000FFF8";
		ram_buffer(3145) := X"24630001";
		ram_buffer(3146) := X"8F828018";
		ram_buffer(3147) := X"03E00008";
		ram_buffer(3148) := X"00000000";
		ram_buffer(3149) := X"8F838038";
		ram_buffer(3150) := X"00000000";
		ram_buffer(3151) := X"10600005";
		ram_buffer(3152) := X"24020001";
		ram_buffer(3153) := X"8F82801C";
		ram_buffer(3154) := X"00000000";
		ram_buffer(3155) := X"2C420001";
		ram_buffer(3156) := X"00021040";
		ram_buffer(3157) := X"03E00008";
		ram_buffer(3158) := X"00000000";
		ram_buffer(3159) := X"1080003E";
		ram_buffer(3160) := X"00000000";
		ram_buffer(3161) := X"8F828018";
		ram_buffer(3162) := X"8C83002C";
		ram_buffer(3163) := X"8C42002C";
		ram_buffer(3164) := X"27BDFFE0";
		ram_buffer(3165) := X"0062102B";
		ram_buffer(3166) := X"AFBF001C";
		ram_buffer(3167) := X"AFB20018";
		ram_buffer(3168) := X"AFB10014";
		ram_buffer(3169) := X"1040002F";
		ram_buffer(3170) := X"AFB00010";
		ram_buffer(3171) := X"8C820018";
		ram_buffer(3172) := X"00000000";
		ram_buffer(3173) := X"04400008";
		ram_buffer(3174) := X"00031080";
		ram_buffer(3175) := X"8F828018";
		ram_buffer(3176) := X"00000000";
		ram_buffer(3177) := X"8C45002C";
		ram_buffer(3178) := X"24020005";
		ram_buffer(3179) := X"00451023";
		ram_buffer(3180) := X"AC820018";
		ram_buffer(3181) := X"00031080";
		ram_buffer(3182) := X"00431021";
		ram_buffer(3183) := X"3C110100";
		ram_buffer(3184) := X"00021080";
		ram_buffer(3185) := X"26315694";
		ram_buffer(3186) := X"8C830014";
		ram_buffer(3187) := X"02221021";
		ram_buffer(3188) := X"14620017";
		ram_buffer(3189) := X"24920004";
		ram_buffer(3190) := X"00808025";
		ram_buffer(3191) := X"0C400545";
		ram_buffer(3192) := X"02402025";
		ram_buffer(3193) := X"8F828018";
		ram_buffer(3194) := X"8F83803C";
		ram_buffer(3195) := X"8C42002C";
		ram_buffer(3196) := X"00000000";
		ram_buffer(3197) := X"0062182B";
		ram_buffer(3198) := X"10600002";
		ram_buffer(3199) := X"AE02002C";
		ram_buffer(3200) := X"AF82803C";
		ram_buffer(3201) := X"00022080";
		ram_buffer(3202) := X"00822021";
		ram_buffer(3203) := X"00042080";
		ram_buffer(3204) := X"8FBF001C";
		ram_buffer(3205) := X"8FB00010";
		ram_buffer(3206) := X"02402825";
		ram_buffer(3207) := X"02242021";
		ram_buffer(3208) := X"8FB20018";
		ram_buffer(3209) := X"8FB10014";
		ram_buffer(3210) := X"0840051C";
		ram_buffer(3211) := X"27BD0020";
		ram_buffer(3212) := X"8F828018";
		ram_buffer(3213) := X"00000000";
		ram_buffer(3214) := X"8C42002C";
		ram_buffer(3215) := X"00000000";
		ram_buffer(3216) := X"AC82002C";
		ram_buffer(3217) := X"8FBF001C";
		ram_buffer(3218) := X"8FB20018";
		ram_buffer(3219) := X"8FB10014";
		ram_buffer(3220) := X"8FB00010";
		ram_buffer(3221) := X"27BD0020";
		ram_buffer(3222) := X"03E00008";
		ram_buffer(3223) := X"00000000";
		ram_buffer(3224) := X"14800009";
		ram_buffer(3225) := X"00001025";
		ram_buffer(3226) := X"03E00008";
		ram_buffer(3227) := X"00000000";
		ram_buffer(3228) := X"00001025";
		ram_buffer(3229) := X"8FBF001C";
		ram_buffer(3230) := X"8FB10018";
		ram_buffer(3231) := X"8FB00014";
		ram_buffer(3232) := X"03E00008";
		ram_buffer(3233) := X"27BD0020";
		ram_buffer(3234) := X"8F828018";
		ram_buffer(3235) := X"27BDFFE0";
		ram_buffer(3236) := X"AFB00014";
		ram_buffer(3237) := X"AFBF001C";
		ram_buffer(3238) := X"AFB10018";
		ram_buffer(3239) := X"10820005";
		ram_buffer(3240) := X"00808025";
		ram_buffer(3241) := X"3C040100";
		ram_buffer(3242) := X"24050ED6";
		ram_buffer(3243) := X"0C40026D";
		ram_buffer(3244) := X"2484552C";
		ram_buffer(3245) := X"8E02004C";
		ram_buffer(3246) := X"00000000";
		ram_buffer(3247) := X"14400005";
		ram_buffer(3248) := X"3C040100";
		ram_buffer(3249) := X"24050ED8";
		ram_buffer(3250) := X"0C40026D";
		ram_buffer(3251) := X"2484552C";
		ram_buffer(3252) := X"8E02004C";
		ram_buffer(3253) := X"8E04002C";
		ram_buffer(3254) := X"8E030048";
		ram_buffer(3255) := X"2442FFFF";
		ram_buffer(3256) := X"1083FFE3";
		ram_buffer(3257) := X"AE02004C";
		ram_buffer(3258) := X"1440FFE2";
		ram_buffer(3259) := X"00001025";
		ram_buffer(3260) := X"26110004";
		ram_buffer(3261) := X"0C400545";
		ram_buffer(3262) := X"02202025";
		ram_buffer(3263) := X"8E040048";
		ram_buffer(3264) := X"24020005";
		ram_buffer(3265) := X"00441023";
		ram_buffer(3266) := X"AE020018";
		ram_buffer(3267) := X"8F82803C";
		ram_buffer(3268) := X"00000000";
		ram_buffer(3269) := X"0044102B";
		ram_buffer(3270) := X"10400002";
		ram_buffer(3271) := X"AE04002C";
		ram_buffer(3272) := X"AF84803C";
		ram_buffer(3273) := X"00041080";
		ram_buffer(3274) := X"00442021";
		ram_buffer(3275) := X"3C020100";
		ram_buffer(3276) := X"24425694";
		ram_buffer(3277) := X"00042080";
		ram_buffer(3278) := X"00442021";
		ram_buffer(3279) := X"0C40051C";
		ram_buffer(3280) := X"02202825";
		ram_buffer(3281) := X"1000FFCB";
		ram_buffer(3282) := X"24020001";
		ram_buffer(3283) := X"27BDFFE8";
		ram_buffer(3284) := X"AFBF0014";
		ram_buffer(3285) := X"0C400284";
		ram_buffer(3286) := X"00000000";
		ram_buffer(3287) := X"8F828038";
		ram_buffer(3288) := X"00000000";
		ram_buffer(3289) := X"10400008";
		ram_buffer(3290) := X"00000000";
		ram_buffer(3291) := X"8F838018";
		ram_buffer(3292) := X"00000000";
		ram_buffer(3293) := X"8C620044";
		ram_buffer(3294) := X"00000000";
		ram_buffer(3295) := X"24420001";
		ram_buffer(3296) := X"AC620044";
		ram_buffer(3297) := X"8F828018";
		ram_buffer(3298) := X"8FBF0014";
		ram_buffer(3299) := X"00000000";
		ram_buffer(3300) := X"03E00008";
		ram_buffer(3301) := X"27BD0018";
		ram_buffer(3302) := X"8F828038";
		ram_buffer(3303) := X"00000000";
		ram_buffer(3304) := X"10400015";
		ram_buffer(3305) := X"00000000";
		ram_buffer(3306) := X"8F828018";
		ram_buffer(3307) := X"00000000";
		ram_buffer(3308) := X"8C420044";
		ram_buffer(3309) := X"00000000";
		ram_buffer(3310) := X"1040000F";
		ram_buffer(3311) := X"00000000";
		ram_buffer(3312) := X"8F838018";
		ram_buffer(3313) := X"00000000";
		ram_buffer(3314) := X"8C620044";
		ram_buffer(3315) := X"00000000";
		ram_buffer(3316) := X"2442FFFF";
		ram_buffer(3317) := X"AC620044";
		ram_buffer(3318) := X"8F828018";
		ram_buffer(3319) := X"00000000";
		ram_buffer(3320) := X"8C420044";
		ram_buffer(3321) := X"00000000";
		ram_buffer(3322) := X"14400003";
		ram_buffer(3323) := X"00000000";
		ram_buffer(3324) := X"0840027F";
		ram_buffer(3325) := X"00000000";
		ram_buffer(3326) := X"03E00008";
		ram_buffer(3327) := X"00000000";
		ram_buffer(3328) := X"27BDFFC8";
		ram_buffer(3329) := X"AFB2001C";
		ram_buffer(3330) := X"00069080";
		ram_buffer(3331) := X"AFB40024";
		ram_buffer(3332) := X"0080A025";
		ram_buffer(3333) := X"02402025";
		ram_buffer(3334) := X"AFB70030";
		ram_buffer(3335) := X"AFB50028";
		ram_buffer(3336) := X"AFB30020";
		ram_buffer(3337) := X"AFB10018";
		ram_buffer(3338) := X"AFBF0034";
		ram_buffer(3339) := X"AFB6002C";
		ram_buffer(3340) := X"AFB00014";
		ram_buffer(3341) := X"00A08825";
		ram_buffer(3342) := X"8FB3004C";
		ram_buffer(3343) := X"0C4012E8";
		ram_buffer(3344) := X"00E0A825";
		ram_buffer(3345) := X"1040008F";
		ram_buffer(3346) := X"2417FFFF";
		ram_buffer(3347) := X"24040058";
		ram_buffer(3348) := X"0C4012E8";
		ram_buffer(3349) := X"0040B025";
		ram_buffer(3350) := X"10400087";
		ram_buffer(3351) := X"00408025";
		ram_buffer(3352) := X"02403025";
		ram_buffer(3353) := X"240500A5";
		ram_buffer(3354) := X"AC560030";
		ram_buffer(3355) := X"0C40146F";
		ram_buffer(3356) := X"02C02025";
		ram_buffer(3357) := X"2642FFFC";
		ram_buffer(3358) := X"8E120030";
		ram_buffer(3359) := X"02202825";
		ram_buffer(3360) := X"02429021";
		ram_buffer(3361) := X"2402FFFC";
		ram_buffer(3362) := X"02429024";
		ram_buffer(3363) := X"26230010";
		ram_buffer(3364) := X"26020034";
		ram_buffer(3365) := X"80A40000";
		ram_buffer(3366) := X"00000000";
		ram_buffer(3367) := X"A0440000";
		ram_buffer(3368) := X"80A40000";
		ram_buffer(3369) := X"00000000";
		ram_buffer(3370) := X"10800003";
		ram_buffer(3371) := X"24A50001";
		ram_buffer(3372) := X"1465FFF8";
		ram_buffer(3373) := X"24420001";
		ram_buffer(3374) := X"8FB60048";
		ram_buffer(3375) := X"00000000";
		ram_buffer(3376) := X"2EC20005";
		ram_buffer(3377) := X"14400002";
		ram_buffer(3378) := X"A2000043";
		ram_buffer(3379) := X"24160004";
		ram_buffer(3380) := X"26110004";
		ram_buffer(3381) := X"AE16002C";
		ram_buffer(3382) := X"AE160048";
		ram_buffer(3383) := X"02202025";
		ram_buffer(3384) := X"0C40051A";
		ram_buffer(3385) := X"AE00004C";
		ram_buffer(3386) := X"0C40051A";
		ram_buffer(3387) := X"26040018";
		ram_buffer(3388) := X"24020005";
		ram_buffer(3389) := X"0056B023";
		ram_buffer(3390) := X"AE000050";
		ram_buffer(3391) := X"AE100010";
		ram_buffer(3392) := X"AE160018";
		ram_buffer(3393) := X"AE100024";
		ram_buffer(3394) := X"AE000044";
		ram_buffer(3395) := X"A2000054";
		ram_buffer(3396) := X"A2000055";
		ram_buffer(3397) := X"02A03025";
		ram_buffer(3398) := X"02802825";
		ram_buffer(3399) := X"0C400085";
		ram_buffer(3400) := X"02402025";
		ram_buffer(3401) := X"12600002";
		ram_buffer(3402) := X"AE020000";
		ram_buffer(3403) := X"AE700000";
		ram_buffer(3404) := X"0C400CD3";
		ram_buffer(3405) := X"00000000";
		ram_buffer(3406) := X"8F828044";
		ram_buffer(3407) := X"3C120100";
		ram_buffer(3408) := X"24420001";
		ram_buffer(3409) := X"AF828044";
		ram_buffer(3410) := X"8F828018";
		ram_buffer(3411) := X"00000000";
		ram_buffer(3412) := X"14400058";
		ram_buffer(3413) := X"00000000";
		ram_buffer(3414) := X"AF908018";
		ram_buffer(3415) := X"8F838044";
		ram_buffer(3416) := X"24020001";
		ram_buffer(3417) := X"14620022";
		ram_buffer(3418) := X"00000000";
		ram_buffer(3419) := X"0C400512";
		ram_buffer(3420) := X"26445694";
		ram_buffer(3421) := X"3C040100";
		ram_buffer(3422) := X"0C400512";
		ram_buffer(3423) := X"248456A8";
		ram_buffer(3424) := X"3C040100";
		ram_buffer(3425) := X"0C400512";
		ram_buffer(3426) := X"248456BC";
		ram_buffer(3427) := X"3C040100";
		ram_buffer(3428) := X"0C400512";
		ram_buffer(3429) := X"248456D0";
		ram_buffer(3430) := X"3C040100";
		ram_buffer(3431) := X"248456E4";
		ram_buffer(3432) := X"0C400512";
		ram_buffer(3433) := X"3C140100";
		ram_buffer(3434) := X"3C130100";
		ram_buffer(3435) := X"0C400512";
		ram_buffer(3436) := X"26845680";
		ram_buffer(3437) := X"0C400512";
		ram_buffer(3438) := X"2664566C";
		ram_buffer(3439) := X"3C040100";
		ram_buffer(3440) := X"0C400512";
		ram_buffer(3441) := X"24845658";
		ram_buffer(3442) := X"3C040100";
		ram_buffer(3443) := X"0C400512";
		ram_buffer(3444) := X"24845644";
		ram_buffer(3445) := X"3C040100";
		ram_buffer(3446) := X"24845630";
		ram_buffer(3447) := X"26945680";
		ram_buffer(3448) := X"0C400512";
		ram_buffer(3449) := X"2673566C";
		ram_buffer(3450) := X"AF948050";
		ram_buffer(3451) := X"AF93804C";
		ram_buffer(3452) := X"8F828028";
		ram_buffer(3453) := X"8E04002C";
		ram_buffer(3454) := X"24420001";
		ram_buffer(3455) := X"AF828028";
		ram_buffer(3456) := X"8F82803C";
		ram_buffer(3457) := X"00000000";
		ram_buffer(3458) := X"0044102B";
		ram_buffer(3459) := X"10400003";
		ram_buffer(3460) := X"00041080";
		ram_buffer(3461) := X"AF84803C";
		ram_buffer(3462) := X"00041080";
		ram_buffer(3463) := X"00441021";
		ram_buffer(3464) := X"00021080";
		ram_buffer(3465) := X"26445694";
		ram_buffer(3466) := X"00822021";
		ram_buffer(3467) := X"0C40051C";
		ram_buffer(3468) := X"02202825";
		ram_buffer(3469) := X"0C400CE6";
		ram_buffer(3470) := X"00000000";
		ram_buffer(3471) := X"8F828038";
		ram_buffer(3472) := X"00000000";
		ram_buffer(3473) := X"1040000F";
		ram_buffer(3474) := X"24170001";
		ram_buffer(3475) := X"8F828018";
		ram_buffer(3476) := X"8E03002C";
		ram_buffer(3477) := X"8C42002C";
		ram_buffer(3478) := X"00000000";
		ram_buffer(3479) := X"0043102B";
		ram_buffer(3480) := X"10400008";
		ram_buffer(3481) := X"00000000";
		ram_buffer(3482) := X"0C400120";
		ram_buffer(3483) := X"00000000";
		ram_buffer(3484) := X"10000004";
		ram_buffer(3485) := X"00000000";
		ram_buffer(3486) := X"0C40135A";
		ram_buffer(3487) := X"02C02025";
		ram_buffer(3488) := X"2417FFFF";
		ram_buffer(3489) := X"8FBF0034";
		ram_buffer(3490) := X"02E01025";
		ram_buffer(3491) := X"8FB6002C";
		ram_buffer(3492) := X"8FB70030";
		ram_buffer(3493) := X"8FB50028";
		ram_buffer(3494) := X"8FB40024";
		ram_buffer(3495) := X"8FB30020";
		ram_buffer(3496) := X"8FB2001C";
		ram_buffer(3497) := X"8FB10018";
		ram_buffer(3498) := X"8FB00014";
		ram_buffer(3499) := X"03E00008";
		ram_buffer(3500) := X"27BD0038";
		ram_buffer(3501) := X"8F828038";
		ram_buffer(3502) := X"00000000";
		ram_buffer(3503) := X"1440FFCC";
		ram_buffer(3504) := X"00000000";
		ram_buffer(3505) := X"8F828018";
		ram_buffer(3506) := X"8E03002C";
		ram_buffer(3507) := X"8C42002C";
		ram_buffer(3508) := X"00000000";
		ram_buffer(3509) := X"0062102B";
		ram_buffer(3510) := X"1440FFC5";
		ram_buffer(3511) := X"00000000";
		ram_buffer(3512) := X"AF908018";
		ram_buffer(3513) := X"1000FFC2";
		ram_buffer(3514) := X"00000000";
		ram_buffer(3515) := X"27BDFFE0";
		ram_buffer(3516) := X"27828020";
		ram_buffer(3517) := X"3C050100";
		ram_buffer(3518) := X"3C040100";
		ram_buffer(3519) := X"00003825";
		ram_buffer(3520) := X"AFA20014";
		ram_buffer(3521) := X"AFA00010";
		ram_buffer(3522) := X"2406012C";
		ram_buffer(3523) := X"24A55544";
		ram_buffer(3524) := X"AFB00018";
		ram_buffer(3525) := X"AFBF001C";
		ram_buffer(3526) := X"0C400D00";
		ram_buffer(3527) := X"248440E4";
		ram_buffer(3528) := X"00408025";
		ram_buffer(3529) := X"24020001";
		ram_buffer(3530) := X"1602000C";
		ram_buffer(3531) := X"2402FFFF";
		ram_buffer(3532) := X"0C400284";
		ram_buffer(3533) := X"00000000";
		ram_buffer(3534) := X"2402FFFF";
		ram_buffer(3535) := X"AF828024";
		ram_buffer(3536) := X"8FBF001C";
		ram_buffer(3537) := X"AF908038";
		ram_buffer(3538) := X"8FB00018";
		ram_buffer(3539) := X"27BD0020";
		ram_buffer(3540) := X"AF808040";
		ram_buffer(3541) := X"084012B4";
		ram_buffer(3542) := X"00000000";
		ram_buffer(3543) := X"16020007";
		ram_buffer(3544) := X"3C040100";
		ram_buffer(3545) := X"8FBF001C";
		ram_buffer(3546) := X"8FB00018";
		ram_buffer(3547) := X"2405078B";
		ram_buffer(3548) := X"2484552C";
		ram_buffer(3549) := X"0840026D";
		ram_buffer(3550) := X"27BD0020";
		ram_buffer(3551) := X"8FBF001C";
		ram_buffer(3552) := X"8FB00018";
		ram_buffer(3553) := X"03E00008";
		ram_buffer(3554) := X"27BD0020";
		ram_buffer(3555) := X"27BDFFE0";
		ram_buffer(3556) := X"AFB00014";
		ram_buffer(3557) := X"00808025";
		ram_buffer(3558) := X"AFBF001C";
		ram_buffer(3559) := X"0C400CD3";
		ram_buffer(3560) := X"AFB10018";
		ram_buffer(3561) := X"16000004";
		ram_buffer(3562) := X"26110004";
		ram_buffer(3563) := X"8F908018";
		ram_buffer(3564) := X"00000000";
		ram_buffer(3565) := X"26110004";
		ram_buffer(3566) := X"0C400545";
		ram_buffer(3567) := X"02202025";
		ram_buffer(3568) := X"8E020028";
		ram_buffer(3569) := X"00000000";
		ram_buffer(3570) := X"10400003";
		ram_buffer(3571) := X"00000000";
		ram_buffer(3572) := X"0C400545";
		ram_buffer(3573) := X"26040018";
		ram_buffer(3574) := X"8F828028";
		ram_buffer(3575) := X"00000000";
		ram_buffer(3576) := X"24420001";
		ram_buffer(3577) := X"AF828028";
		ram_buffer(3578) := X"8F828018";
		ram_buffer(3579) := X"00000000";
		ram_buffer(3580) := X"1602001E";
		ram_buffer(3581) := X"02202825";
		ram_buffer(3582) := X"3C040100";
		ram_buffer(3583) := X"0C40051C";
		ram_buffer(3584) := X"24845644";
		ram_buffer(3585) := X"8F828048";
		ram_buffer(3586) := X"00000000";
		ram_buffer(3587) := X"24420001";
		ram_buffer(3588) := X"AF828048";
		ram_buffer(3589) := X"0C400CE6";
		ram_buffer(3590) := X"00000000";
		ram_buffer(3591) := X"8F828038";
		ram_buffer(3592) := X"00000000";
		ram_buffer(3593) := X"1040001D";
		ram_buffer(3594) := X"00000000";
		ram_buffer(3595) := X"8F828018";
		ram_buffer(3596) := X"00000000";
		ram_buffer(3597) := X"16020019";
		ram_buffer(3598) := X"00000000";
		ram_buffer(3599) := X"8F82801C";
		ram_buffer(3600) := X"00000000";
		ram_buffer(3601) := X"10400004";
		ram_buffer(3602) := X"24050465";
		ram_buffer(3603) := X"3C040100";
		ram_buffer(3604) := X"0C40026D";
		ram_buffer(3605) := X"2484552C";
		ram_buffer(3606) := X"8FBF001C";
		ram_buffer(3607) := X"8FB10018";
		ram_buffer(3608) := X"8FB00014";
		ram_buffer(3609) := X"08400120";
		ram_buffer(3610) := X"27BD0020";
		ram_buffer(3611) := X"8F828044";
		ram_buffer(3612) := X"8E040030";
		ram_buffer(3613) := X"2442FFFF";
		ram_buffer(3614) := X"AF828044";
		ram_buffer(3615) := X"0C40135A";
		ram_buffer(3616) := X"00000000";
		ram_buffer(3617) := X"0C40135A";
		ram_buffer(3618) := X"02002025";
		ram_buffer(3619) := X"0C4009EF";
		ram_buffer(3620) := X"00000000";
		ram_buffer(3621) := X"1000FFDF";
		ram_buffer(3622) := X"00000000";
		ram_buffer(3623) := X"8FBF001C";
		ram_buffer(3624) := X"8FB10018";
		ram_buffer(3625) := X"8FB00014";
		ram_buffer(3626) := X"03E00008";
		ram_buffer(3627) := X"27BD0020";
		ram_buffer(3628) := X"27BDFFE0";
		ram_buffer(3629) := X"AFB10018";
		ram_buffer(3630) := X"AFBF001C";
		ram_buffer(3631) := X"AFB00014";
		ram_buffer(3632) := X"14800005";
		ram_buffer(3633) := X"00808825";
		ram_buffer(3634) := X"3C040100";
		ram_buffer(3635) := X"24050502";
		ram_buffer(3636) := X"0C40026D";
		ram_buffer(3637) := X"2484552C";
		ram_buffer(3638) := X"8F838018";
		ram_buffer(3639) := X"00000000";
		ram_buffer(3640) := X"12230016";
		ram_buffer(3641) := X"00001025";
		ram_buffer(3642) := X"0C400CD3";
		ram_buffer(3643) := X"00000000";
		ram_buffer(3644) := X"8E300014";
		ram_buffer(3645) := X"0C400CE6";
		ram_buffer(3646) := X"00000000";
		ram_buffer(3647) := X"8F838050";
		ram_buffer(3648) := X"00000000";
		ram_buffer(3649) := X"1203000D";
		ram_buffer(3650) := X"24020002";
		ram_buffer(3651) := X"8F83804C";
		ram_buffer(3652) := X"00000000";
		ram_buffer(3653) := X"12030009";
		ram_buffer(3654) := X"00000000";
		ram_buffer(3655) := X"3C020100";
		ram_buffer(3656) := X"24425630";
		ram_buffer(3657) := X"1602000A";
		ram_buffer(3658) := X"3C030100";
		ram_buffer(3659) := X"8E220028";
		ram_buffer(3660) := X"00000000";
		ram_buffer(3661) := X"2C420001";
		ram_buffer(3662) := X"24420002";
		ram_buffer(3663) := X"8FBF001C";
		ram_buffer(3664) := X"8FB10018";
		ram_buffer(3665) := X"8FB00014";
		ram_buffer(3666) := X"03E00008";
		ram_buffer(3667) := X"27BD0020";
		ram_buffer(3668) := X"24635644";
		ram_buffer(3669) := X"1203FFF9";
		ram_buffer(3670) := X"24020004";
		ram_buffer(3671) := X"1200FFF7";
		ram_buffer(3672) := X"00000000";
		ram_buffer(3673) := X"1000FFF5";
		ram_buffer(3674) := X"24020001";
		ram_buffer(3675) := X"27BDFFE8";
		ram_buffer(3676) := X"AFB00010";
		ram_buffer(3677) := X"AFBF0014";
		ram_buffer(3678) := X"0C400CD3";
		ram_buffer(3679) := X"00808025";
		ram_buffer(3680) := X"16000003";
		ram_buffer(3681) := X"02002025";
		ram_buffer(3682) := X"8F848018";
		ram_buffer(3683) := X"00000000";
		ram_buffer(3684) := X"8C90002C";
		ram_buffer(3685) := X"0C400CE6";
		ram_buffer(3686) := X"00000000";
		ram_buffer(3687) := X"8FBF0014";
		ram_buffer(3688) := X"02001025";
		ram_buffer(3689) := X"8FB00010";
		ram_buffer(3690) := X"03E00008";
		ram_buffer(3691) := X"27BD0018";
		ram_buffer(3692) := X"27BDFFD8";
		ram_buffer(3693) := X"2CA20005";
		ram_buffer(3694) := X"AFB2001C";
		ram_buffer(3695) := X"AFB00014";
		ram_buffer(3696) := X"AFBF0024";
		ram_buffer(3697) := X"AFB30020";
		ram_buffer(3698) := X"AFB10018";
		ram_buffer(3699) := X"00808025";
		ram_buffer(3700) := X"14400006";
		ram_buffer(3701) := X"00A09025";
		ram_buffer(3702) := X"3C040100";
		ram_buffer(3703) := X"24050587";
		ram_buffer(3704) := X"0C40026D";
		ram_buffer(3705) := X"2484552C";
		ram_buffer(3706) := X"24120004";
		ram_buffer(3707) := X"0C400CD3";
		ram_buffer(3708) := X"00000000";
		ram_buffer(3709) := X"16000003";
		ram_buffer(3710) := X"00000000";
		ram_buffer(3711) := X"8F908018";
		ram_buffer(3712) := X"00000000";
		ram_buffer(3713) := X"8E020048";
		ram_buffer(3714) := X"00000000";
		ram_buffer(3715) := X"12420035";
		ram_buffer(3716) := X"0052182B";
		ram_buffer(3717) := X"1060003A";
		ram_buffer(3718) := X"00000000";
		ram_buffer(3719) := X"8F838018";
		ram_buffer(3720) := X"00000000";
		ram_buffer(3721) := X"12030007";
		ram_buffer(3722) := X"00008825";
		ram_buffer(3723) := X"8F838018";
		ram_buffer(3724) := X"00000000";
		ram_buffer(3725) := X"8C71002C";
		ram_buffer(3726) := X"00000000";
		ram_buffer(3727) := X"0251882B";
		ram_buffer(3728) := X"3A310001";
		ram_buffer(3729) := X"8E03002C";
		ram_buffer(3730) := X"00000000";
		ram_buffer(3731) := X"14430002";
		ram_buffer(3732) := X"00000000";
		ram_buffer(3733) := X"AE12002C";
		ram_buffer(3734) := X"8E020018";
		ram_buffer(3735) := X"00000000";
		ram_buffer(3736) := X"04400004";
		ram_buffer(3737) := X"AE120048";
		ram_buffer(3738) := X"24050005";
		ram_buffer(3739) := X"00B29023";
		ram_buffer(3740) := X"AE120018";
		ram_buffer(3741) := X"00031080";
		ram_buffer(3742) := X"00431021";
		ram_buffer(3743) := X"3C120100";
		ram_buffer(3744) := X"00021080";
		ram_buffer(3745) := X"26525694";
		ram_buffer(3746) := X"8E030014";
		ram_buffer(3747) := X"02421021";
		ram_buffer(3748) := X"14620010";
		ram_buffer(3749) := X"26130004";
		ram_buffer(3750) := X"0C400545";
		ram_buffer(3751) := X"02602025";
		ram_buffer(3752) := X"8E02002C";
		ram_buffer(3753) := X"8F83803C";
		ram_buffer(3754) := X"00000000";
		ram_buffer(3755) := X"0062182B";
		ram_buffer(3756) := X"10600002";
		ram_buffer(3757) := X"00000000";
		ram_buffer(3758) := X"AF82803C";
		ram_buffer(3759) := X"00022080";
		ram_buffer(3760) := X"00822021";
		ram_buffer(3761) := X"00042080";
		ram_buffer(3762) := X"02602825";
		ram_buffer(3763) := X"0C40051C";
		ram_buffer(3764) := X"02442021";
		ram_buffer(3765) := X"12200003";
		ram_buffer(3766) := X"00000000";
		ram_buffer(3767) := X"0C400120";
		ram_buffer(3768) := X"00000000";
		ram_buffer(3769) := X"8FBF0024";
		ram_buffer(3770) := X"8FB30020";
		ram_buffer(3771) := X"8FB2001C";
		ram_buffer(3772) := X"8FB10018";
		ram_buffer(3773) := X"8FB00014";
		ram_buffer(3774) := X"08400CE6";
		ram_buffer(3775) := X"27BD0028";
		ram_buffer(3776) := X"8F918018";
		ram_buffer(3777) := X"00000000";
		ram_buffer(3778) := X"02118826";
		ram_buffer(3779) := X"1000FFCD";
		ram_buffer(3780) := X"2E310001";
		ram_buffer(3781) := X"27BDFFE0";
		ram_buffer(3782) := X"AFB00014";
		ram_buffer(3783) := X"00808025";
		ram_buffer(3784) := X"AFBF001C";
		ram_buffer(3785) := X"0C400CD3";
		ram_buffer(3786) := X"AFB10018";
		ram_buffer(3787) := X"16000004";
		ram_buffer(3788) := X"26110004";
		ram_buffer(3789) := X"8F908018";
		ram_buffer(3790) := X"00000000";
		ram_buffer(3791) := X"26110004";
		ram_buffer(3792) := X"0C400545";
		ram_buffer(3793) := X"02202025";
		ram_buffer(3794) := X"8E020028";
		ram_buffer(3795) := X"00000000";
		ram_buffer(3796) := X"10400004";
		ram_buffer(3797) := X"02202825";
		ram_buffer(3798) := X"0C400545";
		ram_buffer(3799) := X"26040018";
		ram_buffer(3800) := X"02202825";
		ram_buffer(3801) := X"3C110100";
		ram_buffer(3802) := X"0C40051C";
		ram_buffer(3803) := X"26245630";
		ram_buffer(3804) := X"0C400CE6";
		ram_buffer(3805) := X"00000000";
		ram_buffer(3806) := X"8F828038";
		ram_buffer(3807) := X"00000000";
		ram_buffer(3808) := X"10400007";
		ram_buffer(3809) := X"00000000";
		ram_buffer(3810) := X"0C400CD3";
		ram_buffer(3811) := X"00000000";
		ram_buffer(3812) := X"0C4009EF";
		ram_buffer(3813) := X"00000000";
		ram_buffer(3814) := X"0C400CE6";
		ram_buffer(3815) := X"00000000";
		ram_buffer(3816) := X"8F828018";
		ram_buffer(3817) := X"00000000";
		ram_buffer(3818) := X"16020017";
		ram_buffer(3819) := X"00000000";
		ram_buffer(3820) := X"8F828038";
		ram_buffer(3821) := X"00000000";
		ram_buffer(3822) := X"1040000D";
		ram_buffer(3823) := X"00000000";
		ram_buffer(3824) := X"8F82801C";
		ram_buffer(3825) := X"00000000";
		ram_buffer(3826) := X"10400004";
		ram_buffer(3827) := X"3C040100";
		ram_buffer(3828) := X"2405065E";
		ram_buffer(3829) := X"0C40026D";
		ram_buffer(3830) := X"2484552C";
		ram_buffer(3831) := X"8FBF001C";
		ram_buffer(3832) := X"8FB10018";
		ram_buffer(3833) := X"8FB00014";
		ram_buffer(3834) := X"08400120";
		ram_buffer(3835) := X"27BD0020";
		ram_buffer(3836) := X"8F828044";
		ram_buffer(3837) := X"8E235630";
		ram_buffer(3838) := X"00000000";
		ram_buffer(3839) := X"14620007";
		ram_buffer(3840) := X"00000000";
		ram_buffer(3841) := X"AF808018";
		ram_buffer(3842) := X"8FBF001C";
		ram_buffer(3843) := X"8FB10018";
		ram_buffer(3844) := X"8FB00014";
		ram_buffer(3845) := X"03E00008";
		ram_buffer(3846) := X"27BD0020";
		ram_buffer(3847) := X"8FBF001C";
		ram_buffer(3848) := X"8FB10018";
		ram_buffer(3849) := X"8FB00014";
		ram_buffer(3850) := X"08400B3F";
		ram_buffer(3851) := X"27BD0020";
		ram_buffer(3852) := X"14800029";
		ram_buffer(3853) := X"240506B2";
		ram_buffer(3854) := X"3C040100";
		ram_buffer(3855) := X"0840026D";
		ram_buffer(3856) := X"2484552C";
		ram_buffer(3857) := X"0C400CD3";
		ram_buffer(3858) := X"00808025";
		ram_buffer(3859) := X"0C400A02";
		ram_buffer(3860) := X"02002025";
		ram_buffer(3861) := X"1040001B";
		ram_buffer(3862) := X"26110004";
		ram_buffer(3863) := X"0C400545";
		ram_buffer(3864) := X"02202025";
		ram_buffer(3865) := X"8E04002C";
		ram_buffer(3866) := X"8F82803C";
		ram_buffer(3867) := X"00000000";
		ram_buffer(3868) := X"0044102B";
		ram_buffer(3869) := X"10400003";
		ram_buffer(3870) := X"00041080";
		ram_buffer(3871) := X"AF84803C";
		ram_buffer(3872) := X"00041080";
		ram_buffer(3873) := X"00441021";
		ram_buffer(3874) := X"3C040100";
		ram_buffer(3875) := X"00021080";
		ram_buffer(3876) := X"24845694";
		ram_buffer(3877) := X"00822021";
		ram_buffer(3878) := X"0C40051C";
		ram_buffer(3879) := X"02202825";
		ram_buffer(3880) := X"8F838018";
		ram_buffer(3881) := X"8E02002C";
		ram_buffer(3882) := X"8C63002C";
		ram_buffer(3883) := X"00000000";
		ram_buffer(3884) := X"0043102B";
		ram_buffer(3885) := X"14400003";
		ram_buffer(3886) := X"00000000";
		ram_buffer(3887) := X"0C400120";
		ram_buffer(3888) := X"00000000";
		ram_buffer(3889) := X"8FBF001C";
		ram_buffer(3890) := X"8FB10018";
		ram_buffer(3891) := X"8FB00014";
		ram_buffer(3892) := X"08400CE6";
		ram_buffer(3893) := X"27BD0020";
		ram_buffer(3894) := X"8F828018";
		ram_buffer(3895) := X"27BDFFE0";
		ram_buffer(3896) := X"AFBF001C";
		ram_buffer(3897) := X"AFB10018";
		ram_buffer(3898) := X"1482FFD6";
		ram_buffer(3899) := X"AFB00014";
		ram_buffer(3900) := X"8FBF001C";
		ram_buffer(3901) := X"8FB10018";
		ram_buffer(3902) := X"8FB00014";
		ram_buffer(3903) := X"03E00008";
		ram_buffer(3904) := X"27BD0020";
		ram_buffer(3905) := X"8F82801C";
		ram_buffer(3906) := X"27BDFFD0";
		ram_buffer(3907) := X"AFBF002C";
		ram_buffer(3908) := X"AFB50028";
		ram_buffer(3909) := X"AFB40024";
		ram_buffer(3910) := X"AFB30020";
		ram_buffer(3911) := X"AFB2001C";
		ram_buffer(3912) := X"AFB10018";
		ram_buffer(3913) := X"14400005";
		ram_buffer(3914) := X"AFB00014";
		ram_buffer(3915) := X"3C040100";
		ram_buffer(3916) := X"240507EF";
		ram_buffer(3917) := X"0C40026D";
		ram_buffer(3918) := X"2484552C";
		ram_buffer(3919) := X"0C400CD3";
		ram_buffer(3920) := X"00000000";
		ram_buffer(3921) := X"8F82801C";
		ram_buffer(3922) := X"00000000";
		ram_buffer(3923) := X"2442FFFF";
		ram_buffer(3924) := X"AF82801C";
		ram_buffer(3925) := X"8F82801C";
		ram_buffer(3926) := X"00000000";
		ram_buffer(3927) := X"1040000E";
		ram_buffer(3928) := X"00000000";
		ram_buffer(3929) := X"00008025";
		ram_buffer(3930) := X"0C400CE6";
		ram_buffer(3931) := X"00000000";
		ram_buffer(3932) := X"8FBF002C";
		ram_buffer(3933) := X"02001025";
		ram_buffer(3934) := X"8FB50028";
		ram_buffer(3935) := X"8FB40024";
		ram_buffer(3936) := X"8FB30020";
		ram_buffer(3937) := X"8FB2001C";
		ram_buffer(3938) := X"8FB10018";
		ram_buffer(3939) := X"8FB00014";
		ram_buffer(3940) := X"03E00008";
		ram_buffer(3941) := X"27BD0030";
		ram_buffer(3942) := X"8F828044";
		ram_buffer(3943) := X"00000000";
		ram_buffer(3944) := X"1040FFF0";
		ram_buffer(3945) := X"3C140100";
		ram_buffer(3946) := X"3C110100";
		ram_buffer(3947) := X"00008025";
		ram_buffer(3948) := X"26925658";
		ram_buffer(3949) := X"26315694";
		ram_buffer(3950) := X"24130001";
		ram_buffer(3951) := X"8E825658";
		ram_buffer(3952) := X"00000000";
		ram_buffer(3953) := X"1440001A";
		ram_buffer(3954) := X"00000000";
		ram_buffer(3955) := X"12000003";
		ram_buffer(3956) := X"00000000";
		ram_buffer(3957) := X"0C4009EF";
		ram_buffer(3958) := X"00000000";
		ram_buffer(3959) := X"8F908034";
		ram_buffer(3960) := X"00000000";
		ram_buffer(3961) := X"1200000A";
		ram_buffer(3962) := X"24110001";
		ram_buffer(3963) := X"0C400AC4";
		ram_buffer(3964) := X"00000000";
		ram_buffer(3965) := X"10400002";
		ram_buffer(3966) := X"00000000";
		ram_buffer(3967) := X"AF918030";
		ram_buffer(3968) := X"2610FFFF";
		ram_buffer(3969) := X"1600FFF9";
		ram_buffer(3970) := X"00000000";
		ram_buffer(3971) := X"AF808034";
		ram_buffer(3972) := X"8F828030";
		ram_buffer(3973) := X"00000000";
		ram_buffer(3974) := X"1040FFD2";
		ram_buffer(3975) := X"00000000";
		ram_buffer(3976) := X"0C400120";
		ram_buffer(3977) := X"24100001";
		ram_buffer(3978) := X"1000FFCF";
		ram_buffer(3979) := X"00000000";
		ram_buffer(3980) := X"8E42000C";
		ram_buffer(3981) := X"00000000";
		ram_buffer(3982) := X"8C50000C";
		ram_buffer(3983) := X"00000000";
		ram_buffer(3984) := X"26040018";
		ram_buffer(3985) := X"0C400545";
		ram_buffer(3986) := X"26150004";
		ram_buffer(3987) := X"0C400545";
		ram_buffer(3988) := X"02A02025";
		ram_buffer(3989) := X"8E02002C";
		ram_buffer(3990) := X"8F83803C";
		ram_buffer(3991) := X"00000000";
		ram_buffer(3992) := X"0062182B";
		ram_buffer(3993) := X"10600002";
		ram_buffer(3994) := X"00000000";
		ram_buffer(3995) := X"AF82803C";
		ram_buffer(3996) := X"00022080";
		ram_buffer(3997) := X"00822021";
		ram_buffer(3998) := X"00042080";
		ram_buffer(3999) := X"02A02825";
		ram_buffer(4000) := X"0C40051C";
		ram_buffer(4001) := X"02242021";
		ram_buffer(4002) := X"8F838018";
		ram_buffer(4003) := X"8E02002C";
		ram_buffer(4004) := X"8C63002C";
		ram_buffer(4005) := X"00000000";
		ram_buffer(4006) := X"0043102B";
		ram_buffer(4007) := X"1440FFC7";
		ram_buffer(4008) := X"00000000";
		ram_buffer(4009) := X"AF938030";
		ram_buffer(4010) := X"1000FFC4";
		ram_buffer(4011) := X"00000000";
		ram_buffer(4012) := X"27BDFFE0";
		ram_buffer(4013) := X"AFB10018";
		ram_buffer(4014) := X"AFB00014";
		ram_buffer(4015) := X"AFBF001C";
		ram_buffer(4016) := X"00808825";
		ram_buffer(4017) := X"14800005";
		ram_buffer(4018) := X"00A08025";
		ram_buffer(4019) := X"3C040100";
		ram_buffer(4020) := X"24050479";
		ram_buffer(4021) := X"0C40026D";
		ram_buffer(4022) := X"2484552C";
		ram_buffer(4023) := X"16000004";
		ram_buffer(4024) := X"2405047A";
		ram_buffer(4025) := X"3C040100";
		ram_buffer(4026) := X"0C40026D";
		ram_buffer(4027) := X"2484552C";
		ram_buffer(4028) := X"8F82801C";
		ram_buffer(4029) := X"00000000";
		ram_buffer(4030) := X"10400004";
		ram_buffer(4031) := X"3C040100";
		ram_buffer(4032) := X"2405047B";
		ram_buffer(4033) := X"0C40026D";
		ram_buffer(4034) := X"2484552C";
		ram_buffer(4035) := X"0C400A98";
		ram_buffer(4036) := X"00000000";
		ram_buffer(4037) := X"8E230000";
		ram_buffer(4038) := X"8F848040";
		ram_buffer(4039) := X"02038021";
		ram_buffer(4040) := X"0083282B";
		ram_buffer(4041) := X"10A00005";
		ram_buffer(4042) := X"0203182B";
		ram_buffer(4043) := X"10600005";
		ram_buffer(4044) := X"00002825";
		ram_buffer(4045) := X"10000003";
		ram_buffer(4046) := X"0090282B";
		ram_buffer(4047) := X"1060FFFD";
		ram_buffer(4048) := X"24050001";
		ram_buffer(4049) := X"10A00004";
		ram_buffer(4050) := X"AE300000";
		ram_buffer(4051) := X"00002825";
		ram_buffer(4052) := X"0C400A1A";
		ram_buffer(4053) := X"02042023";
		ram_buffer(4054) := X"0C400F41";
		ram_buffer(4055) := X"00000000";
		ram_buffer(4056) := X"14400006";
		ram_buffer(4057) := X"00000000";
		ram_buffer(4058) := X"8FBF001C";
		ram_buffer(4059) := X"8FB10018";
		ram_buffer(4060) := X"8FB00014";
		ram_buffer(4061) := X"08400120";
		ram_buffer(4062) := X"27BD0020";
		ram_buffer(4063) := X"8FBF001C";
		ram_buffer(4064) := X"8FB10018";
		ram_buffer(4065) := X"8FB00014";
		ram_buffer(4066) := X"03E00008";
		ram_buffer(4067) := X"27BD0020";
		ram_buffer(4068) := X"14800007";
		ram_buffer(4069) := X"00000000";
		ram_buffer(4070) := X"08400120";
		ram_buffer(4071) := X"00000000";
		ram_buffer(4072) := X"8FBF0014";
		ram_buffer(4073) := X"8FB00010";
		ram_buffer(4074) := X"1000FFFB";
		ram_buffer(4075) := X"27BD0018";
		ram_buffer(4076) := X"8F82801C";
		ram_buffer(4077) := X"27BDFFE8";
		ram_buffer(4078) := X"AFB00010";
		ram_buffer(4079) := X"AFBF0014";
		ram_buffer(4080) := X"10400005";
		ram_buffer(4081) := X"00808025";
		ram_buffer(4082) := X"3C040100";
		ram_buffer(4083) := X"240504D6";
		ram_buffer(4084) := X"0C40026D";
		ram_buffer(4085) := X"2484552C";
		ram_buffer(4086) := X"0C400A98";
		ram_buffer(4087) := X"00002825";
		ram_buffer(4088) := X"0C400A1A";
		ram_buffer(4089) := X"02002025";
		ram_buffer(4090) := X"0C400F41";
		ram_buffer(4091) := X"00000000";
		ram_buffer(4092) := X"1040FFEB";
		ram_buffer(4093) := X"00000000";
		ram_buffer(4094) := X"8FBF0014";
		ram_buffer(4095) := X"8FB00010";
		ram_buffer(4096) := X"03E00008";
		ram_buffer(4097) := X"27BD0018";
		ram_buffer(4098) := X"27BDFFE0";
		ram_buffer(4099) := X"AFB10018";
		ram_buffer(4100) := X"AFBF001C";
		ram_buffer(4101) := X"AFB00014";
		ram_buffer(4102) := X"0C4014B6";
		ram_buffer(4103) := X"00808825";
		ram_buffer(4104) := X"2C420010";
		ram_buffer(4105) := X"14400004";
		ram_buffer(4106) := X"240508DD";
		ram_buffer(4107) := X"3C040100";
		ram_buffer(4108) := X"0C40026D";
		ram_buffer(4109) := X"2484552C";
		ram_buffer(4110) := X"0C400A98";
		ram_buffer(4111) := X"3C0D0100";
		ram_buffer(4112) := X"00006025";
		ram_buffer(4113) := X"25AD5694";
		ram_buffer(4114) := X"240EFF9C";
		ram_buffer(4115) := X"25840050";
		ram_buffer(4116) := X"02202825";
		ram_buffer(4117) := X"0C4009C2";
		ram_buffer(4118) := X"01A42021";
		ram_buffer(4119) := X"14400019";
		ram_buffer(4120) := X"00408025";
		ram_buffer(4121) := X"258CFFEC";
		ram_buffer(4122) := X"158EFFF9";
		ram_buffer(4123) := X"25840050";
		ram_buffer(4124) := X"8F848050";
		ram_buffer(4125) := X"0C4009C2";
		ram_buffer(4126) := X"02202825";
		ram_buffer(4127) := X"14400011";
		ram_buffer(4128) := X"00408025";
		ram_buffer(4129) := X"8F84804C";
		ram_buffer(4130) := X"0C4009C2";
		ram_buffer(4131) := X"02202825";
		ram_buffer(4132) := X"1440000C";
		ram_buffer(4133) := X"00408025";
		ram_buffer(4134) := X"3C040100";
		ram_buffer(4135) := X"02202825";
		ram_buffer(4136) := X"0C4009C2";
		ram_buffer(4137) := X"24845630";
		ram_buffer(4138) := X"14400006";
		ram_buffer(4139) := X"00408025";
		ram_buffer(4140) := X"3C040100";
		ram_buffer(4141) := X"02202825";
		ram_buffer(4142) := X"0C4009C2";
		ram_buffer(4143) := X"24845644";
		ram_buffer(4144) := X"00408025";
		ram_buffer(4145) := X"0C400F41";
		ram_buffer(4146) := X"00000000";
		ram_buffer(4147) := X"8FBF001C";
		ram_buffer(4148) := X"02001025";
		ram_buffer(4149) := X"8FB10018";
		ram_buffer(4150) := X"8FB00014";
		ram_buffer(4151) := X"03E00008";
		ram_buffer(4152) := X"27BD0020";
		ram_buffer(4153) := X"27BDFFD8";
		ram_buffer(4154) := X"AFB10018";
		ram_buffer(4155) := X"3C110100";
		ram_buffer(4156) := X"AFB30020";
		ram_buffer(4157) := X"AFB2001C";
		ram_buffer(4158) := X"AFBF0024";
		ram_buffer(4159) := X"AFB00014";
		ram_buffer(4160) := X"26335644";
		ram_buffer(4161) := X"3C120100";
		ram_buffer(4162) := X"8F828048";
		ram_buffer(4163) := X"00000000";
		ram_buffer(4164) := X"1440000A";
		ram_buffer(4165) := X"00000000";
		ram_buffer(4166) := X"8E425694";
		ram_buffer(4167) := X"00000000";
		ram_buffer(4168) := X"2C420002";
		ram_buffer(4169) := X"1440FFF8";
		ram_buffer(4170) := X"00000000";
		ram_buffer(4171) := X"0C400120";
		ram_buffer(4172) := X"00000000";
		ram_buffer(4173) := X"1000FFF4";
		ram_buffer(4174) := X"00000000";
		ram_buffer(4175) := X"0C400A98";
		ram_buffer(4176) := X"00000000";
		ram_buffer(4177) := X"8E305644";
		ram_buffer(4178) := X"0C400F41";
		ram_buffer(4179) := X"00000000";
		ram_buffer(4180) := X"1200FFED";
		ram_buffer(4181) := X"00000000";
		ram_buffer(4182) := X"0C400CD3";
		ram_buffer(4183) := X"00000000";
		ram_buffer(4184) := X"8E62000C";
		ram_buffer(4185) := X"00000000";
		ram_buffer(4186) := X"8C50000C";
		ram_buffer(4187) := X"0C400545";
		ram_buffer(4188) := X"26040004";
		ram_buffer(4189) := X"8F828044";
		ram_buffer(4190) := X"00000000";
		ram_buffer(4191) := X"2442FFFF";
		ram_buffer(4192) := X"AF828044";
		ram_buffer(4193) := X"8F828048";
		ram_buffer(4194) := X"00000000";
		ram_buffer(4195) := X"2442FFFF";
		ram_buffer(4196) := X"AF828048";
		ram_buffer(4197) := X"0C400CE6";
		ram_buffer(4198) := X"00000000";
		ram_buffer(4199) := X"8E040030";
		ram_buffer(4200) := X"0C40135A";
		ram_buffer(4201) := X"00000000";
		ram_buffer(4202) := X"0C40135A";
		ram_buffer(4203) := X"02002025";
		ram_buffer(4204) := X"1000FFD5";
		ram_buffer(4205) := X"00000000";
		ram_buffer(4206) := X"27BDFFE0";
		ram_buffer(4207) := X"AFB00014";
		ram_buffer(4208) := X"AFBF001C";
		ram_buffer(4209) := X"AFB10018";
		ram_buffer(4210) := X"14800005";
		ram_buffer(4211) := X"00808025";
		ram_buffer(4212) := X"3C040100";
		ram_buffer(4213) := X"24050987";
		ram_buffer(4214) := X"0C40026D";
		ram_buffer(4215) := X"2484552C";
		ram_buffer(4216) := X"0C400A98";
		ram_buffer(4217) := X"02002025";
		ram_buffer(4218) := X"0C400E2C";
		ram_buffer(4219) := X"00000000";
		ram_buffer(4220) := X"24030002";
		ram_buffer(4221) := X"14430026";
		ram_buffer(4222) := X"26110004";
		ram_buffer(4223) := X"0C400545";
		ram_buffer(4224) := X"02202025";
		ram_buffer(4225) := X"0C400CD3";
		ram_buffer(4226) := X"00000000";
		ram_buffer(4227) := X"8E020028";
		ram_buffer(4228) := X"00000000";
		ram_buffer(4229) := X"10400005";
		ram_buffer(4230) := X"00000000";
		ram_buffer(4231) := X"0C400545";
		ram_buffer(4232) := X"26040018";
		ram_buffer(4233) := X"24020001";
		ram_buffer(4234) := X"A2020055";
		ram_buffer(4235) := X"0C400CE6";
		ram_buffer(4236) := X"00000000";
		ram_buffer(4237) := X"8E04002C";
		ram_buffer(4238) := X"8F82803C";
		ram_buffer(4239) := X"00000000";
		ram_buffer(4240) := X"0044102B";
		ram_buffer(4241) := X"10400003";
		ram_buffer(4242) := X"00041080";
		ram_buffer(4243) := X"AF84803C";
		ram_buffer(4244) := X"00041080";
		ram_buffer(4245) := X"00441021";
		ram_buffer(4246) := X"3C040100";
		ram_buffer(4247) := X"00021080";
		ram_buffer(4248) := X"24845694";
		ram_buffer(4249) := X"00822021";
		ram_buffer(4250) := X"0C40051C";
		ram_buffer(4251) := X"02202825";
		ram_buffer(4252) := X"8F838018";
		ram_buffer(4253) := X"8E02002C";
		ram_buffer(4254) := X"8C63002C";
		ram_buffer(4255) := X"00000000";
		ram_buffer(4256) := X"0062102B";
		ram_buffer(4257) := X"10400002";
		ram_buffer(4258) := X"24020001";
		ram_buffer(4259) := X"AF828030";
		ram_buffer(4260) := X"0C400F41";
		ram_buffer(4261) := X"00000000";
		ram_buffer(4262) := X"8FBF001C";
		ram_buffer(4263) := X"8FB10018";
		ram_buffer(4264) := X"8FB00014";
		ram_buffer(4265) := X"00001025";
		ram_buffer(4266) := X"03E00008";
		ram_buffer(4267) := X"27BD0020";
		ram_buffer(4268) := X"27BDFFE0";
		ram_buffer(4269) := X"AFB20018";
		ram_buffer(4270) := X"AFB10014";
		ram_buffer(4271) := X"AFBF001C";
		ram_buffer(4272) := X"AFB00010";
		ram_buffer(4273) := X"00808825";
		ram_buffer(4274) := X"14800005";
		ram_buffer(4275) := X"00A09025";
		ram_buffer(4276) := X"3C040100";
		ram_buffer(4277) := X"24050BDA";
		ram_buffer(4278) := X"0C40026D";
		ram_buffer(4279) := X"2484552C";
		ram_buffer(4280) := X"16400004";
		ram_buffer(4281) := X"3C040100";
		ram_buffer(4282) := X"24050BDB";
		ram_buffer(4283) := X"0C40026D";
		ram_buffer(4284) := X"2484552C";
		ram_buffer(4285) := X"0C400CD3";
		ram_buffer(4286) := X"00000000";
		ram_buffer(4287) := X"8F848040";
		ram_buffer(4288) := X"8F828018";
		ram_buffer(4289) := X"00000000";
		ram_buffer(4290) := X"90420055";
		ram_buffer(4291) := X"00000000";
		ram_buffer(4292) := X"1040000D";
		ram_buffer(4293) := X"2402FFFF";
		ram_buffer(4294) := X"8F828018";
		ram_buffer(4295) := X"24100001";
		ram_buffer(4296) := X"A0400055";
		ram_buffer(4297) := X"0C400CE6";
		ram_buffer(4298) := X"00000000";
		ram_buffer(4299) := X"8FBF001C";
		ram_buffer(4300) := X"02001025";
		ram_buffer(4301) := X"8FB20018";
		ram_buffer(4302) := X"8FB10014";
		ram_buffer(4303) := X"8FB00010";
		ram_buffer(4304) := X"03E00008";
		ram_buffer(4305) := X"27BD0020";
		ram_buffer(4306) := X"8E430000";
		ram_buffer(4307) := X"00000000";
		ram_buffer(4308) := X"1062FFF4";
		ram_buffer(4309) := X"00008025";
		ram_buffer(4310) := X"8F85802C";
		ram_buffer(4311) := X"8E260000";
		ram_buffer(4312) := X"8E220004";
		ram_buffer(4313) := X"10C50003";
		ram_buffer(4314) := X"0082282B";
		ram_buffer(4315) := X"10A0FFED";
		ram_buffer(4316) := X"24100001";
		ram_buffer(4317) := X"00822823";
		ram_buffer(4318) := X"00A3282B";
		ram_buffer(4319) := X"10A0FFE9";
		ram_buffer(4320) := X"24100001";
		ram_buffer(4321) := X"00641823";
		ram_buffer(4322) := X"00621821";
		ram_buffer(4323) := X"AE430000";
		ram_buffer(4324) := X"0C400C24";
		ram_buffer(4325) := X"02202025";
		ram_buffer(4326) := X"1000FFE2";
		ram_buffer(4327) := X"00008025";
		ram_buffer(4328) := X"8F828018";
		ram_buffer(4329) := X"8F848018";
		ram_buffer(4330) := X"8F838018";
		ram_buffer(4331) := X"8C420018";
		ram_buffer(4332) := X"8C65002C";
		ram_buffer(4333) := X"24030005";
		ram_buffer(4334) := X"00651823";
		ram_buffer(4335) := X"03E00008";
		ram_buffer(4336) := X"AC830018";
		ram_buffer(4337) := X"8F828018";
		ram_buffer(4338) := X"00000000";
		ram_buffer(4339) := X"10400007";
		ram_buffer(4340) := X"00000000";
		ram_buffer(4341) := X"8F838018";
		ram_buffer(4342) := X"00000000";
		ram_buffer(4343) := X"8C62004C";
		ram_buffer(4344) := X"00000000";
		ram_buffer(4345) := X"24420001";
		ram_buffer(4346) := X"AC62004C";
		ram_buffer(4347) := X"8F828018";
		ram_buffer(4348) := X"03E00008";
		ram_buffer(4349) := X"00000000";
		ram_buffer(4350) := X"27BDFFE0";
		ram_buffer(4351) := X"AFB10018";
		ram_buffer(4352) := X"AFB00014";
		ram_buffer(4353) := X"AFBF001C";
		ram_buffer(4354) := X"00808825";
		ram_buffer(4355) := X"0C400CD3";
		ram_buffer(4356) := X"00A08025";
		ram_buffer(4357) := X"8F828018";
		ram_buffer(4358) := X"00000000";
		ram_buffer(4359) := X"8C420050";
		ram_buffer(4360) := X"00000000";
		ram_buffer(4361) := X"1440000A";
		ram_buffer(4362) := X"00000000";
		ram_buffer(4363) := X"8F828018";
		ram_buffer(4364) := X"24030001";
		ram_buffer(4365) := X"A0430054";
		ram_buffer(4366) := X"12000005";
		ram_buffer(4367) := X"24050001";
		ram_buffer(4368) := X"0C400A1A";
		ram_buffer(4369) := X"02002025";
		ram_buffer(4370) := X"0C400120";
		ram_buffer(4371) := X"00000000";
		ram_buffer(4372) := X"0C400CE6";
		ram_buffer(4373) := X"00000000";
		ram_buffer(4374) := X"0C400CD3";
		ram_buffer(4375) := X"00000000";
		ram_buffer(4376) := X"8F828018";
		ram_buffer(4377) := X"00000000";
		ram_buffer(4378) := X"8C500050";
		ram_buffer(4379) := X"00000000";
		ram_buffer(4380) := X"12000005";
		ram_buffer(4381) := X"00000000";
		ram_buffer(4382) := X"8F828018";
		ram_buffer(4383) := X"1220000D";
		ram_buffer(4384) := X"2603FFFF";
		ram_buffer(4385) := X"AC400050";
		ram_buffer(4386) := X"8F828018";
		ram_buffer(4387) := X"00000000";
		ram_buffer(4388) := X"A0400054";
		ram_buffer(4389) := X"0C400CE6";
		ram_buffer(4390) := X"00000000";
		ram_buffer(4391) := X"8FBF001C";
		ram_buffer(4392) := X"02001025";
		ram_buffer(4393) := X"8FB10018";
		ram_buffer(4394) := X"8FB00014";
		ram_buffer(4395) := X"03E00008";
		ram_buffer(4396) := X"27BD0020";
		ram_buffer(4397) := X"AC430050";
		ram_buffer(4398) := X"1000FFF3";
		ram_buffer(4399) := X"00000000";
		ram_buffer(4400) := X"27BDFFD8";
		ram_buffer(4401) := X"AFB30020";
		ram_buffer(4402) := X"AFB2001C";
		ram_buffer(4403) := X"AFB10018";
		ram_buffer(4404) := X"AFB00014";
		ram_buffer(4405) := X"AFBF0024";
		ram_buffer(4406) := X"00808825";
		ram_buffer(4407) := X"00A08025";
		ram_buffer(4408) := X"00C09025";
		ram_buffer(4409) := X"0C400CD3";
		ram_buffer(4410) := X"00E09825";
		ram_buffer(4411) := X"8F828018";
		ram_buffer(4412) := X"24030002";
		ram_buffer(4413) := X"90420054";
		ram_buffer(4414) := X"00000000";
		ram_buffer(4415) := X"304200FF";
		ram_buffer(4416) := X"10430010";
		ram_buffer(4417) := X"00000000";
		ram_buffer(4418) := X"8F828018";
		ram_buffer(4419) := X"00118827";
		ram_buffer(4420) := X"8C440050";
		ram_buffer(4421) := X"24030001";
		ram_buffer(4422) := X"02248824";
		ram_buffer(4423) := X"AC510050";
		ram_buffer(4424) := X"8F828018";
		ram_buffer(4425) := X"00000000";
		ram_buffer(4426) := X"A0430054";
		ram_buffer(4427) := X"12600005";
		ram_buffer(4428) := X"24050001";
		ram_buffer(4429) := X"0C400A1A";
		ram_buffer(4430) := X"02602025";
		ram_buffer(4431) := X"0C400120";
		ram_buffer(4432) := X"00000000";
		ram_buffer(4433) := X"0C400CE6";
		ram_buffer(4434) := X"00000000";
		ram_buffer(4435) := X"0C400CD3";
		ram_buffer(4436) := X"00000000";
		ram_buffer(4437) := X"12400006";
		ram_buffer(4438) := X"00000000";
		ram_buffer(4439) := X"8F828018";
		ram_buffer(4440) := X"00000000";
		ram_buffer(4441) := X"8C420050";
		ram_buffer(4442) := X"00000000";
		ram_buffer(4443) := X"AE420000";
		ram_buffer(4444) := X"8F828018";
		ram_buffer(4445) := X"00008825";
		ram_buffer(4446) := X"90430054";
		ram_buffer(4447) := X"24020001";
		ram_buffer(4448) := X"306300FF";
		ram_buffer(4449) := X"10620007";
		ram_buffer(4450) := X"00000000";
		ram_buffer(4451) := X"8F828018";
		ram_buffer(4452) := X"00108027";
		ram_buffer(4453) := X"8C430050";
		ram_buffer(4454) := X"24110001";
		ram_buffer(4455) := X"02038024";
		ram_buffer(4456) := X"AC500050";
		ram_buffer(4457) := X"8F828018";
		ram_buffer(4458) := X"00000000";
		ram_buffer(4459) := X"A0400054";
		ram_buffer(4460) := X"0C400CE6";
		ram_buffer(4461) := X"00000000";
		ram_buffer(4462) := X"8FBF0024";
		ram_buffer(4463) := X"02201025";
		ram_buffer(4464) := X"8FB30020";
		ram_buffer(4465) := X"8FB2001C";
		ram_buffer(4466) := X"8FB10018";
		ram_buffer(4467) := X"8FB00014";
		ram_buffer(4468) := X"03E00008";
		ram_buffer(4469) := X"27BD0028";
		ram_buffer(4470) := X"27BDFFD8";
		ram_buffer(4471) := X"AFB30020";
		ram_buffer(4472) := X"AFB2001C";
		ram_buffer(4473) := X"AFB10018";
		ram_buffer(4474) := X"AFB00014";
		ram_buffer(4475) := X"AFBF0024";
		ram_buffer(4476) := X"00808025";
		ram_buffer(4477) := X"00A09025";
		ram_buffer(4478) := X"00C08825";
		ram_buffer(4479) := X"14800005";
		ram_buffer(4480) := X"00E09825";
		ram_buffer(4481) := X"3C040100";
		ram_buffer(4482) := X"2405110C";
		ram_buffer(4483) := X"0C40026D";
		ram_buffer(4484) := X"2484552C";
		ram_buffer(4485) := X"0C400CD3";
		ram_buffer(4486) := X"00000000";
		ram_buffer(4487) := X"12600004";
		ram_buffer(4488) := X"00000000";
		ram_buffer(4489) := X"8E020050";
		ram_buffer(4490) := X"00000000";
		ram_buffer(4491) := X"AE620000";
		ram_buffer(4492) := X"92030054";
		ram_buffer(4493) := X"24020002";
		ram_buffer(4494) := X"A2020054";
		ram_buffer(4495) := X"24020002";
		ram_buffer(4496) := X"12220023";
		ram_buffer(4497) := X"306300FF";
		ram_buffer(4498) := X"2E240003";
		ram_buffer(4499) := X"10800009";
		ram_buffer(4500) := X"00000000";
		ram_buffer(4501) := X"24020001";
		ram_buffer(4502) := X"12220017";
		ram_buffer(4503) := X"00000000";
		ram_buffer(4504) := X"24020001";
		ram_buffer(4505) := X"10620020";
		ram_buffer(4506) := X"00000000";
		ram_buffer(4507) := X"10000008";
		ram_buffer(4508) := X"24110001";
		ram_buffer(4509) := X"24040003";
		ram_buffer(4510) := X"12240012";
		ram_buffer(4511) := X"24040004";
		ram_buffer(4512) := X"1624FFF7";
		ram_buffer(4513) := X"00000000";
		ram_buffer(4514) := X"1462000E";
		ram_buffer(4515) := X"00008825";
		ram_buffer(4516) := X"0C400CE6";
		ram_buffer(4517) := X"00000000";
		ram_buffer(4518) := X"8FBF0024";
		ram_buffer(4519) := X"02201025";
		ram_buffer(4520) := X"8FB30020";
		ram_buffer(4521) := X"8FB2001C";
		ram_buffer(4522) := X"8FB10018";
		ram_buffer(4523) := X"8FB00014";
		ram_buffer(4524) := X"03E00008";
		ram_buffer(4525) := X"27BD0028";
		ram_buffer(4526) := X"8E020050";
		ram_buffer(4527) := X"00000000";
		ram_buffer(4528) := X"00529025";
		ram_buffer(4529) := X"AE120050";
		ram_buffer(4530) := X"1000FFE6";
		ram_buffer(4531) := X"24020001";
		ram_buffer(4532) := X"8E020050";
		ram_buffer(4533) := X"00000000";
		ram_buffer(4534) := X"24420001";
		ram_buffer(4535) := X"AE020050";
		ram_buffer(4536) := X"1000FFE0";
		ram_buffer(4537) := X"24020001";
		ram_buffer(4538) := X"26110004";
		ram_buffer(4539) := X"0C400545";
		ram_buffer(4540) := X"02202025";
		ram_buffer(4541) := X"8E04002C";
		ram_buffer(4542) := X"8F82803C";
		ram_buffer(4543) := X"00000000";
		ram_buffer(4544) := X"0044102B";
		ram_buffer(4545) := X"10400003";
		ram_buffer(4546) := X"00041080";
		ram_buffer(4547) := X"AF84803C";
		ram_buffer(4548) := X"00041080";
		ram_buffer(4549) := X"00441021";
		ram_buffer(4550) := X"3C040100";
		ram_buffer(4551) := X"00021080";
		ram_buffer(4552) := X"24845694";
		ram_buffer(4553) := X"00822021";
		ram_buffer(4554) := X"0C40051C";
		ram_buffer(4555) := X"02202825";
		ram_buffer(4556) := X"8E020028";
		ram_buffer(4557) := X"00000000";
		ram_buffer(4558) := X"10400004";
		ram_buffer(4559) := X"3C040100";
		ram_buffer(4560) := X"24051144";
		ram_buffer(4561) := X"0C40026D";
		ram_buffer(4562) := X"2484552C";
		ram_buffer(4563) := X"8F838018";
		ram_buffer(4564) := X"8E02002C";
		ram_buffer(4565) := X"8C63002C";
		ram_buffer(4566) := X"00000000";
		ram_buffer(4567) := X"0062102B";
		ram_buffer(4568) := X"1040FFC2";
		ram_buffer(4569) := X"00000000";
		ram_buffer(4570) := X"0C400120";
		ram_buffer(4571) := X"24110001";
		ram_buffer(4572) := X"1000FFC7";
		ram_buffer(4573) := X"00000000";
		ram_buffer(4574) := X"27BDFFD8";
		ram_buffer(4575) := X"AFB40020";
		ram_buffer(4576) := X"AFB3001C";
		ram_buffer(4577) := X"AFB20018";
		ram_buffer(4578) := X"AFB10014";
		ram_buffer(4579) := X"AFB00010";
		ram_buffer(4580) := X"AFBF0024";
		ram_buffer(4581) := X"00808025";
		ram_buffer(4582) := X"00A09825";
		ram_buffer(4583) := X"00C08825";
		ram_buffer(4584) := X"8FB20038";
		ram_buffer(4585) := X"14800005";
		ram_buffer(4586) := X"00E0A025";
		ram_buffer(4587) := X"3C040100";
		ram_buffer(4588) := X"24051177";
		ram_buffer(4589) := X"0C40026D";
		ram_buffer(4590) := X"2484552C";
		ram_buffer(4591) := X"12800004";
		ram_buffer(4592) := X"00000000";
		ram_buffer(4593) := X"8E020050";
		ram_buffer(4594) := X"00000000";
		ram_buffer(4595) := X"AE820000";
		ram_buffer(4596) := X"92030054";
		ram_buffer(4597) := X"24020002";
		ram_buffer(4598) := X"24040002";
		ram_buffer(4599) := X"306300FF";
		ram_buffer(4600) := X"A2020054";
		ram_buffer(4601) := X"12240021";
		ram_buffer(4602) := X"00000000";
		ram_buffer(4603) := X"2E220003";
		ram_buffer(4604) := X"10400009";
		ram_buffer(4605) := X"24020003";
		ram_buffer(4606) := X"24020001";
		ram_buffer(4607) := X"12220015";
		ram_buffer(4608) := X"00000000";
		ram_buffer(4609) := X"24020001";
		ram_buffer(4610) := X"1062001E";
		ram_buffer(4611) := X"00000000";
		ram_buffer(4612) := X"10000008";
		ram_buffer(4613) := X"24020001";
		ram_buffer(4614) := X"12220011";
		ram_buffer(4615) := X"00000000";
		ram_buffer(4616) := X"24020004";
		ram_buffer(4617) := X"1622FFF7";
		ram_buffer(4618) := X"00000000";
		ram_buffer(4619) := X"1464000C";
		ram_buffer(4620) := X"00001025";
		ram_buffer(4621) := X"8FBF0024";
		ram_buffer(4622) := X"8FB40020";
		ram_buffer(4623) := X"8FB3001C";
		ram_buffer(4624) := X"8FB20018";
		ram_buffer(4625) := X"8FB10014";
		ram_buffer(4626) := X"8FB00010";
		ram_buffer(4627) := X"03E00008";
		ram_buffer(4628) := X"27BD0028";
		ram_buffer(4629) := X"8E020050";
		ram_buffer(4630) := X"00000000";
		ram_buffer(4631) := X"00539825";
		ram_buffer(4632) := X"AE130050";
		ram_buffer(4633) := X"1000FFE8";
		ram_buffer(4634) := X"24020001";
		ram_buffer(4635) := X"8E020050";
		ram_buffer(4636) := X"00000000";
		ram_buffer(4637) := X"24420001";
		ram_buffer(4638) := X"AE020050";
		ram_buffer(4639) := X"1000FFE2";
		ram_buffer(4640) := X"24020001";
		ram_buffer(4641) := X"8E020028";
		ram_buffer(4642) := X"00000000";
		ram_buffer(4643) := X"10400004";
		ram_buffer(4644) := X"240511BE";
		ram_buffer(4645) := X"3C040100";
		ram_buffer(4646) := X"0C40026D";
		ram_buffer(4647) := X"2484552C";
		ram_buffer(4648) := X"8F82801C";
		ram_buffer(4649) := X"00000000";
		ram_buffer(4650) := X"1440001F";
		ram_buffer(4651) := X"3C040100";
		ram_buffer(4652) := X"26110004";
		ram_buffer(4653) := X"0C400545";
		ram_buffer(4654) := X"02202025";
		ram_buffer(4655) := X"8E04002C";
		ram_buffer(4656) := X"8F82803C";
		ram_buffer(4657) := X"00000000";
		ram_buffer(4658) := X"0044102B";
		ram_buffer(4659) := X"10400003";
		ram_buffer(4660) := X"00041080";
		ram_buffer(4661) := X"AF84803C";
		ram_buffer(4662) := X"00041080";
		ram_buffer(4663) := X"00441021";
		ram_buffer(4664) := X"3C040100";
		ram_buffer(4665) := X"00021080";
		ram_buffer(4666) := X"24845694";
		ram_buffer(4667) := X"02202825";
		ram_buffer(4668) := X"00822021";
		ram_buffer(4669) := X"0C40051C";
		ram_buffer(4670) := X"00000000";
		ram_buffer(4671) := X"8F838018";
		ram_buffer(4672) := X"8E02002C";
		ram_buffer(4673) := X"8C63002C";
		ram_buffer(4674) := X"00000000";
		ram_buffer(4675) := X"0062102B";
		ram_buffer(4676) := X"1040FFBF";
		ram_buffer(4677) := X"00000000";
		ram_buffer(4678) := X"12400006";
		ram_buffer(4679) := X"24020001";
		ram_buffer(4680) := X"1000FFC4";
		ram_buffer(4681) := X"AE420000";
		ram_buffer(4682) := X"26050018";
		ram_buffer(4683) := X"1000FFF1";
		ram_buffer(4684) := X"24845658";
		ram_buffer(4685) := X"AF828030";
		ram_buffer(4686) := X"1000FFBE";
		ram_buffer(4687) := X"00000000";
		ram_buffer(4688) := X"27BDFFE0";
		ram_buffer(4689) := X"AFB10014";
		ram_buffer(4690) := X"AFB00010";
		ram_buffer(4691) := X"AFBF001C";
		ram_buffer(4692) := X"AFB20018";
		ram_buffer(4693) := X"00808025";
		ram_buffer(4694) := X"14800005";
		ram_buffer(4695) := X"00A08825";
		ram_buffer(4696) := X"3C040100";
		ram_buffer(4697) := X"240511F2";
		ram_buffer(4698) := X"0C40026D";
		ram_buffer(4699) := X"2484552C";
		ram_buffer(4700) := X"24030002";
		ram_buffer(4701) := X"92020054";
		ram_buffer(4702) := X"A2030054";
		ram_buffer(4703) := X"8E030050";
		ram_buffer(4704) := X"304200FF";
		ram_buffer(4705) := X"24630001";
		ram_buffer(4706) := X"AE030050";
		ram_buffer(4707) := X"24030001";
		ram_buffer(4708) := X"14430029";
		ram_buffer(4709) := X"00000000";
		ram_buffer(4710) := X"8E020028";
		ram_buffer(4711) := X"00000000";
		ram_buffer(4712) := X"10400004";
		ram_buffer(4713) := X"24051218";
		ram_buffer(4714) := X"3C040100";
		ram_buffer(4715) := X"0C40026D";
		ram_buffer(4716) := X"2484552C";
		ram_buffer(4717) := X"8F82801C";
		ram_buffer(4718) := X"00000000";
		ram_buffer(4719) := X"14400024";
		ram_buffer(4720) := X"3C040100";
		ram_buffer(4721) := X"26120004";
		ram_buffer(4722) := X"0C400545";
		ram_buffer(4723) := X"02402025";
		ram_buffer(4724) := X"8E04002C";
		ram_buffer(4725) := X"8F82803C";
		ram_buffer(4726) := X"00000000";
		ram_buffer(4727) := X"0044102B";
		ram_buffer(4728) := X"10400003";
		ram_buffer(4729) := X"00041080";
		ram_buffer(4730) := X"AF84803C";
		ram_buffer(4731) := X"00041080";
		ram_buffer(4732) := X"00441021";
		ram_buffer(4733) := X"3C040100";
		ram_buffer(4734) := X"00021080";
		ram_buffer(4735) := X"24845694";
		ram_buffer(4736) := X"02402825";
		ram_buffer(4737) := X"00822021";
		ram_buffer(4738) := X"0C40051C";
		ram_buffer(4739) := X"00000000";
		ram_buffer(4740) := X"8F838018";
		ram_buffer(4741) := X"8E02002C";
		ram_buffer(4742) := X"8C63002C";
		ram_buffer(4743) := X"00000000";
		ram_buffer(4744) := X"0062102B";
		ram_buffer(4745) := X"10400004";
		ram_buffer(4746) := X"00000000";
		ram_buffer(4747) := X"1220000B";
		ram_buffer(4748) := X"24020001";
		ram_buffer(4749) := X"AE220000";
		ram_buffer(4750) := X"8FBF001C";
		ram_buffer(4751) := X"8FB20018";
		ram_buffer(4752) := X"8FB10014";
		ram_buffer(4753) := X"8FB00010";
		ram_buffer(4754) := X"03E00008";
		ram_buffer(4755) := X"27BD0020";
		ram_buffer(4756) := X"26050018";
		ram_buffer(4757) := X"1000FFEC";
		ram_buffer(4758) := X"24845658";
		ram_buffer(4759) := X"AF828030";
		ram_buffer(4760) := X"1000FFF5";
		ram_buffer(4761) := X"00000000";
		ram_buffer(4762) := X"27BDFFE0";
		ram_buffer(4763) := X"AFB00014";
		ram_buffer(4764) := X"AFBF001C";
		ram_buffer(4765) := X"AFB10018";
		ram_buffer(4766) := X"14800002";
		ram_buffer(4767) := X"00808025";
		ram_buffer(4768) := X"8F908018";
		ram_buffer(4769) := X"0C400CD3";
		ram_buffer(4770) := X"00000000";
		ram_buffer(4771) := X"92030054";
		ram_buffer(4772) := X"24020002";
		ram_buffer(4773) := X"306300FF";
		ram_buffer(4774) := X"14620003";
		ram_buffer(4775) := X"00008825";
		ram_buffer(4776) := X"A2000054";
		ram_buffer(4777) := X"24110001";
		ram_buffer(4778) := X"0C400CE6";
		ram_buffer(4779) := X"00000000";
		ram_buffer(4780) := X"8FBF001C";
		ram_buffer(4781) := X"02201025";
		ram_buffer(4782) := X"8FB00014";
		ram_buffer(4783) := X"8FB10018";
		ram_buffer(4784) := X"03E00008";
		ram_buffer(4785) := X"27BD0020";
		ram_buffer(4786) := X"03E00008";
		ram_buffer(4787) := X"00000000";
		ram_buffer(4788) := X"27BDFFE8";
		ram_buffer(4789) := X"AFBF0014";
		ram_buffer(4790) := X"0C4000E7";
		ram_buffer(4791) := X"00000000";
		ram_buffer(4792) := X"0C40027F";
		ram_buffer(4793) := X"00000000";
		ram_buffer(4794) := X"0C4000F6";
		ram_buffer(4795) := X"00000000";
		ram_buffer(4796) := X"0C400284";
		ram_buffer(4797) := X"00000000";
		ram_buffer(4798) := X"1000FFFF";
		ram_buffer(4799) := X"00000000";
		ram_buffer(4800) := X"3C040100";
		ram_buffer(4801) := X"24050070";
		ram_buffer(4802) := X"0840026D";
		ram_buffer(4803) := X"2484554C";
		ram_buffer(4804) := X"27828068";
		ram_buffer(4805) := X"8C430000";
		ram_buffer(4806) := X"00000000";
		ram_buffer(4807) := X"0064282B";
		ram_buffer(4808) := X"14A0001D";
		ram_buffer(4809) := X"00000000";
		ram_buffer(4810) := X"8C450004";
		ram_buffer(4811) := X"00000000";
		ram_buffer(4812) := X"00453021";
		ram_buffer(4813) := X"14860006";
		ram_buffer(4814) := X"00000000";
		ram_buffer(4815) := X"8C840004";
		ram_buffer(4816) := X"00000000";
		ram_buffer(4817) := X"00852021";
		ram_buffer(4818) := X"AC440004";
		ram_buffer(4819) := X"00402025";
		ram_buffer(4820) := X"8C860004";
		ram_buffer(4821) := X"00000000";
		ram_buffer(4822) := X"00862821";
		ram_buffer(4823) := X"14650009";
		ram_buffer(4824) := X"00000000";
		ram_buffer(4825) := X"8F858064";
		ram_buffer(4826) := X"00000000";
		ram_buffer(4827) := X"10650005";
		ram_buffer(4828) := X"00000000";
		ram_buffer(4829) := X"8C650004";
		ram_buffer(4830) := X"8C630000";
		ram_buffer(4831) := X"00A62821";
		ram_buffer(4832) := X"AC850004";
		ram_buffer(4833) := X"10820002";
		ram_buffer(4834) := X"AC830000";
		ram_buffer(4835) := X"AC440000";
		ram_buffer(4836) := X"03E00008";
		ram_buffer(4837) := X"00000000";
		ram_buffer(4838) := X"1000FFDE";
		ram_buffer(4839) := X"00601025";
		ram_buffer(4840) := X"27BDFFD8";
		ram_buffer(4841) := X"AFB00014";
		ram_buffer(4842) := X"AFBF0024";
		ram_buffer(4843) := X"AFB30020";
		ram_buffer(4844) := X"AFB2001C";
		ram_buffer(4845) := X"AFB10018";
		ram_buffer(4846) := X"0C400A98";
		ram_buffer(4847) := X"00808025";
		ram_buffer(4848) := X"8F828064";
		ram_buffer(4849) := X"00000000";
		ram_buffer(4850) := X"14400012";
		ram_buffer(4851) := X"3C050100";
		ram_buffer(4852) := X"24A356F8";
		ram_buffer(4853) := X"3402FFF8";
		ram_buffer(4854) := X"2404FFFC";
		ram_buffer(4855) := X"00621021";
		ram_buffer(4856) := X"00441024";
		ram_buffer(4857) := X"00432023";
		ram_buffer(4858) := X"AF80806C";
		ram_buffer(4859) := X"AF838068";
		ram_buffer(4860) := X"AC400004";
		ram_buffer(4861) := X"AC400000";
		ram_buffer(4862) := X"AF828064";
		ram_buffer(4863) := X"ACA256F8";
		ram_buffer(4864) := X"3C028000";
		ram_buffer(4865) := X"AC640004";
		ram_buffer(4866) := X"AF84805C";
		ram_buffer(4867) := X"AF848060";
		ram_buffer(4868) := X"AF828058";
		ram_buffer(4869) := X"8F828058";
		ram_buffer(4870) := X"00000000";
		ram_buffer(4871) := X"02021024";
		ram_buffer(4872) := X"1440003A";
		ram_buffer(4873) := X"00009025";
		ram_buffer(4874) := X"12000038";
		ram_buffer(4875) := X"26100008";
		ram_buffer(4876) := X"32020003";
		ram_buffer(4877) := X"10400003";
		ram_buffer(4878) := X"2404FFFC";
		ram_buffer(4879) := X"02048024";
		ram_buffer(4880) := X"26100004";
		ram_buffer(4881) := X"12000031";
		ram_buffer(4882) := X"00009025";
		ram_buffer(4883) := X"8F828060";
		ram_buffer(4884) := X"00000000";
		ram_buffer(4885) := X"0050102B";
		ram_buffer(4886) := X"1440002C";
		ram_buffer(4887) := X"27838068";
		ram_buffer(4888) := X"8F918068";
		ram_buffer(4889) := X"00000000";
		ram_buffer(4890) := X"8E220004";
		ram_buffer(4891) := X"00000000";
		ram_buffer(4892) := X"0050202B";
		ram_buffer(4893) := X"14800035";
		ram_buffer(4894) := X"00000000";
		ram_buffer(4895) := X"8F848064";
		ram_buffer(4896) := X"00000000";
		ram_buffer(4897) := X"12240021";
		ram_buffer(4898) := X"00009025";
		ram_buffer(4899) := X"8C720000";
		ram_buffer(4900) := X"8E240000";
		ram_buffer(4901) := X"00501023";
		ram_buffer(4902) := X"2C420011";
		ram_buffer(4903) := X"26520008";
		ram_buffer(4904) := X"1440000E";
		ram_buffer(4905) := X"AC640000";
		ram_buffer(4906) := X"02309821";
		ram_buffer(4907) := X"32620003";
		ram_buffer(4908) := X"10400004";
		ram_buffer(4909) := X"3C040100";
		ram_buffer(4910) := X"240500EC";
		ram_buffer(4911) := X"0C40026D";
		ram_buffer(4912) := X"24845564";
		ram_buffer(4913) := X"8E220004";
		ram_buffer(4914) := X"02602025";
		ram_buffer(4915) := X"00501023";
		ram_buffer(4916) := X"AE620004";
		ram_buffer(4917) := X"0C4012C4";
		ram_buffer(4918) := X"AE300004";
		ram_buffer(4919) := X"8F828060";
		ram_buffer(4920) := X"8E240004";
		ram_buffer(4921) := X"8F83805C";
		ram_buffer(4922) := X"00441023";
		ram_buffer(4923) := X"0043182B";
		ram_buffer(4924) := X"10600002";
		ram_buffer(4925) := X"AF828060";
		ram_buffer(4926) := X"AF82805C";
		ram_buffer(4927) := X"8F828058";
		ram_buffer(4928) := X"AE200000";
		ram_buffer(4929) := X"00441025";
		ram_buffer(4930) := X"AE220004";
		ram_buffer(4931) := X"0C400F41";
		ram_buffer(4932) := X"00000000";
		ram_buffer(4933) := X"32420003";
		ram_buffer(4934) := X"10400004";
		ram_buffer(4935) := X"2405012C";
		ram_buffer(4936) := X"3C040100";
		ram_buffer(4937) := X"0C40026D";
		ram_buffer(4938) := X"24845564";
		ram_buffer(4939) := X"8FBF0024";
		ram_buffer(4940) := X"02401025";
		ram_buffer(4941) := X"8FB30020";
		ram_buffer(4942) := X"8FB2001C";
		ram_buffer(4943) := X"8FB10018";
		ram_buffer(4944) := X"8FB00014";
		ram_buffer(4945) := X"03E00008";
		ram_buffer(4946) := X"27BD0028";
		ram_buffer(4947) := X"8E240000";
		ram_buffer(4948) := X"00000000";
		ram_buffer(4949) := X"1080FFC9";
		ram_buffer(4950) := X"00000000";
		ram_buffer(4951) := X"02201825";
		ram_buffer(4952) := X"1000FFC1";
		ram_buffer(4953) := X"00808825";
		ram_buffer(4954) := X"1080002E";
		ram_buffer(4955) := X"00000000";
		ram_buffer(4956) := X"8C82FFFC";
		ram_buffer(4957) := X"8F838058";
		ram_buffer(4958) := X"27BDFFE8";
		ram_buffer(4959) := X"00431024";
		ram_buffer(4960) := X"AFB00010";
		ram_buffer(4961) := X"AFBF0014";
		ram_buffer(4962) := X"14400005";
		ram_buffer(4963) := X"00808025";
		ram_buffer(4964) := X"3C040100";
		ram_buffer(4965) := X"24050140";
		ram_buffer(4966) := X"0C40026D";
		ram_buffer(4967) := X"24845564";
		ram_buffer(4968) := X"8E02FFF8";
		ram_buffer(4969) := X"00000000";
		ram_buffer(4970) := X"10400004";
		ram_buffer(4971) := X"3C040100";
		ram_buffer(4972) := X"24050141";
		ram_buffer(4973) := X"0C40026D";
		ram_buffer(4974) := X"24845564";
		ram_buffer(4975) := X"8E03FFFC";
		ram_buffer(4976) := X"8F828058";
		ram_buffer(4977) := X"00000000";
		ram_buffer(4978) := X"00622024";
		ram_buffer(4979) := X"10800012";
		ram_buffer(4980) := X"00000000";
		ram_buffer(4981) := X"8E04FFF8";
		ram_buffer(4982) := X"00000000";
		ram_buffer(4983) := X"1480000E";
		ram_buffer(4984) := X"00021027";
		ram_buffer(4985) := X"00431024";
		ram_buffer(4986) := X"0C400A98";
		ram_buffer(4987) := X"AE02FFFC";
		ram_buffer(4988) := X"8E03FFFC";
		ram_buffer(4989) := X"8F828060";
		ram_buffer(4990) := X"2604FFF8";
		ram_buffer(4991) := X"00431021";
		ram_buffer(4992) := X"0C4012C4";
		ram_buffer(4993) := X"AF828060";
		ram_buffer(4994) := X"8FBF0014";
		ram_buffer(4995) := X"8FB00010";
		ram_buffer(4996) := X"08400F41";
		ram_buffer(4997) := X"27BD0018";
		ram_buffer(4998) := X"8FBF0014";
		ram_buffer(4999) := X"8FB00010";
		ram_buffer(5000) := X"27BD0018";
		ram_buffer(5001) := X"03E00008";
		ram_buffer(5002) := X"00000000";
		ram_buffer(5003) := X"8F828060";
		ram_buffer(5004) := X"03E00008";
		ram_buffer(5005) := X"00000000";
		ram_buffer(5006) := X"8F82805C";
		ram_buffer(5007) := X"03E00008";
		ram_buffer(5008) := X"00000000";
		ram_buffer(5009) := X"03E00008";
		ram_buffer(5010) := X"00000000";
		ram_buffer(5011) := X"28CA0008";
		ram_buffer(5012) := X"1540005B";
		ram_buffer(5013) := X"00801025";
		ram_buffer(5014) := X"00A4C026";
		ram_buffer(5015) := X"33180003";
		ram_buffer(5016) := X"17000066";
		ram_buffer(5017) := X"00043823";
		ram_buffer(5018) := X"30E70003";
		ram_buffer(5019) := X"10E00005";
		ram_buffer(5020) := X"00C73023";
		ram_buffer(5021) := X"88B80000";
		ram_buffer(5022) := X"00A72821";
		ram_buffer(5023) := X"A8980000";
		ram_buffer(5024) := X"00872021";
		ram_buffer(5025) := X"30D8003F";
		ram_buffer(5026) := X"10D80026";
		ram_buffer(5027) := X"00D83823";
		ram_buffer(5028) := X"00873821";
		ram_buffer(5029) := X"8CA80000";
		ram_buffer(5030) := X"8CA90004";
		ram_buffer(5031) := X"8CAA0008";
		ram_buffer(5032) := X"8CAB000C";
		ram_buffer(5033) := X"8CAC0010";
		ram_buffer(5034) := X"8CAD0014";
		ram_buffer(5035) := X"8CAE0018";
		ram_buffer(5036) := X"8CAF001C";
		ram_buffer(5037) := X"AC880000";
		ram_buffer(5038) := X"AC890004";
		ram_buffer(5039) := X"AC8A0008";
		ram_buffer(5040) := X"AC8B000C";
		ram_buffer(5041) := X"AC8C0010";
		ram_buffer(5042) := X"AC8D0014";
		ram_buffer(5043) := X"AC8E0018";
		ram_buffer(5044) := X"AC8F001C";
		ram_buffer(5045) := X"8CA80020";
		ram_buffer(5046) := X"8CA90024";
		ram_buffer(5047) := X"8CAA0028";
		ram_buffer(5048) := X"8CAB002C";
		ram_buffer(5049) := X"8CAC0030";
		ram_buffer(5050) := X"8CAD0034";
		ram_buffer(5051) := X"8CAE0038";
		ram_buffer(5052) := X"8CAF003C";
		ram_buffer(5053) := X"AC880020";
		ram_buffer(5054) := X"AC890024";
		ram_buffer(5055) := X"AC8A0028";
		ram_buffer(5056) := X"AC8B002C";
		ram_buffer(5057) := X"AC8C0030";
		ram_buffer(5058) := X"AC8D0034";
		ram_buffer(5059) := X"AC8E0038";
		ram_buffer(5060) := X"AC8F003C";
		ram_buffer(5061) := X"24840040";
		ram_buffer(5062) := X"1487FFDE";
		ram_buffer(5063) := X"24A50040";
		ram_buffer(5064) := X"03003025";
		ram_buffer(5065) := X"30D8001F";
		ram_buffer(5066) := X"10D80013";
		ram_buffer(5067) := X"00000000";
		ram_buffer(5068) := X"8CA80000";
		ram_buffer(5069) := X"8CA90004";
		ram_buffer(5070) := X"8CAA0008";
		ram_buffer(5071) := X"8CAB000C";
		ram_buffer(5072) := X"8CAC0010";
		ram_buffer(5073) := X"8CAD0014";
		ram_buffer(5074) := X"8CAE0018";
		ram_buffer(5075) := X"8CAF001C";
		ram_buffer(5076) := X"24A50020";
		ram_buffer(5077) := X"AC880000";
		ram_buffer(5078) := X"AC890004";
		ram_buffer(5079) := X"AC8A0008";
		ram_buffer(5080) := X"AC8B000C";
		ram_buffer(5081) := X"AC8C0010";
		ram_buffer(5082) := X"AC8D0014";
		ram_buffer(5083) := X"AC8E0018";
		ram_buffer(5084) := X"AC8F001C";
		ram_buffer(5085) := X"24840020";
		ram_buffer(5086) := X"33060003";
		ram_buffer(5087) := X"10D80007";
		ram_buffer(5088) := X"03063823";
		ram_buffer(5089) := X"00873821";
		ram_buffer(5090) := X"8CAB0000";
		ram_buffer(5091) := X"24840004";
		ram_buffer(5092) := X"24A50004";
		ram_buffer(5093) := X"1487FFFC";
		ram_buffer(5094) := X"AC8BFFFC";
		ram_buffer(5095) := X"18C00006";
		ram_buffer(5096) := X"00863821";
		ram_buffer(5097) := X"80A30000";
		ram_buffer(5098) := X"24840001";
		ram_buffer(5099) := X"24A50001";
		ram_buffer(5100) := X"1487FFFC";
		ram_buffer(5101) := X"A083FFFF";
		ram_buffer(5102) := X"03E00008";
		ram_buffer(5103) := X"00000000";
		ram_buffer(5104) := X"30D80003";
		ram_buffer(5105) := X"1306FFF5";
		ram_buffer(5106) := X"30990003";
		ram_buffer(5107) := X"1720FFF3";
		ram_buffer(5108) := X"30B90003";
		ram_buffer(5109) := X"1720FFF1";
		ram_buffer(5110) := X"00D83823";
		ram_buffer(5111) := X"00873821";
		ram_buffer(5112) := X"8CAB0000";
		ram_buffer(5113) := X"24840004";
		ram_buffer(5114) := X"24A50004";
		ram_buffer(5115) := X"1487FFFC";
		ram_buffer(5116) := X"AC8BFFFC";
		ram_buffer(5117) := X"1000FFE9";
		ram_buffer(5118) := X"03003025";
		ram_buffer(5119) := X"30E70003";
		ram_buffer(5120) := X"10E00006";
		ram_buffer(5121) := X"00C73023";
		ram_buffer(5122) := X"88A30000";
		ram_buffer(5123) := X"98A30003";
		ram_buffer(5124) := X"00A72821";
		ram_buffer(5125) := X"A8830000";
		ram_buffer(5126) := X"00872021";
		ram_buffer(5127) := X"30D8003F";
		ram_buffer(5128) := X"10D80036";
		ram_buffer(5129) := X"00D83823";
		ram_buffer(5130) := X"00873821";
		ram_buffer(5131) := X"88A80000";
		ram_buffer(5132) := X"88A90004";
		ram_buffer(5133) := X"88AA0008";
		ram_buffer(5134) := X"88AB000C";
		ram_buffer(5135) := X"88AC0010";
		ram_buffer(5136) := X"88AD0014";
		ram_buffer(5137) := X"88AE0018";
		ram_buffer(5138) := X"88AF001C";
		ram_buffer(5139) := X"98A80003";
		ram_buffer(5140) := X"98A90007";
		ram_buffer(5141) := X"98AA000B";
		ram_buffer(5142) := X"98AB000F";
		ram_buffer(5143) := X"98AC0013";
		ram_buffer(5144) := X"98AD0017";
		ram_buffer(5145) := X"98AE001B";
		ram_buffer(5146) := X"98AF001F";
		ram_buffer(5147) := X"AC880000";
		ram_buffer(5148) := X"AC890004";
		ram_buffer(5149) := X"AC8A0008";
		ram_buffer(5150) := X"AC8B000C";
		ram_buffer(5151) := X"AC8C0010";
		ram_buffer(5152) := X"AC8D0014";
		ram_buffer(5153) := X"AC8E0018";
		ram_buffer(5154) := X"AC8F001C";
		ram_buffer(5155) := X"88A80020";
		ram_buffer(5156) := X"88A90024";
		ram_buffer(5157) := X"88AA0028";
		ram_buffer(5158) := X"88AB002C";
		ram_buffer(5159) := X"88AC0030";
		ram_buffer(5160) := X"88AD0034";
		ram_buffer(5161) := X"88AE0038";
		ram_buffer(5162) := X"88AF003C";
		ram_buffer(5163) := X"98A80023";
		ram_buffer(5164) := X"98A90027";
		ram_buffer(5165) := X"98AA002B";
		ram_buffer(5166) := X"98AB002F";
		ram_buffer(5167) := X"98AC0033";
		ram_buffer(5168) := X"98AD0037";
		ram_buffer(5169) := X"98AE003B";
		ram_buffer(5170) := X"98AF003F";
		ram_buffer(5171) := X"AC880020";
		ram_buffer(5172) := X"AC890024";
		ram_buffer(5173) := X"AC8A0028";
		ram_buffer(5174) := X"AC8B002C";
		ram_buffer(5175) := X"AC8C0030";
		ram_buffer(5176) := X"AC8D0034";
		ram_buffer(5177) := X"AC8E0038";
		ram_buffer(5178) := X"AC8F003C";
		ram_buffer(5179) := X"24840040";
		ram_buffer(5180) := X"1487FFCE";
		ram_buffer(5181) := X"24A50040";
		ram_buffer(5182) := X"03003025";
		ram_buffer(5183) := X"30D8001F";
		ram_buffer(5184) := X"10D8001B";
		ram_buffer(5185) := X"00000000";
		ram_buffer(5186) := X"88A80000";
		ram_buffer(5187) := X"88A90004";
		ram_buffer(5188) := X"88AA0008";
		ram_buffer(5189) := X"88AB000C";
		ram_buffer(5190) := X"88AC0010";
		ram_buffer(5191) := X"88AD0014";
		ram_buffer(5192) := X"88AE0018";
		ram_buffer(5193) := X"88AF001C";
		ram_buffer(5194) := X"98A80003";
		ram_buffer(5195) := X"98A90007";
		ram_buffer(5196) := X"98AA000B";
		ram_buffer(5197) := X"98AB000F";
		ram_buffer(5198) := X"98AC0013";
		ram_buffer(5199) := X"98AD0017";
		ram_buffer(5200) := X"98AE001B";
		ram_buffer(5201) := X"98AF001F";
		ram_buffer(5202) := X"24A50020";
		ram_buffer(5203) := X"AC880000";
		ram_buffer(5204) := X"AC890004";
		ram_buffer(5205) := X"AC8A0008";
		ram_buffer(5206) := X"AC8B000C";
		ram_buffer(5207) := X"AC8C0010";
		ram_buffer(5208) := X"AC8D0014";
		ram_buffer(5209) := X"AC8E0018";
		ram_buffer(5210) := X"AC8F001C";
		ram_buffer(5211) := X"24840020";
		ram_buffer(5212) := X"33060003";
		ram_buffer(5213) := X"10D80008";
		ram_buffer(5214) := X"03063823";
		ram_buffer(5215) := X"00873821";
		ram_buffer(5216) := X"88A30000";
		ram_buffer(5217) := X"98A30003";
		ram_buffer(5218) := X"24840004";
		ram_buffer(5219) := X"24A50004";
		ram_buffer(5220) := X"1487FFFB";
		ram_buffer(5221) := X"AC83FFFC";
		ram_buffer(5222) := X"10C0FF87";
		ram_buffer(5223) := X"00863821";
		ram_buffer(5224) := X"80A30000";
		ram_buffer(5225) := X"24840001";
		ram_buffer(5226) := X"24A50001";
		ram_buffer(5227) := X"1487FFFC";
		ram_buffer(5228) := X"A083FFFF";
		ram_buffer(5229) := X"03E00008";
		ram_buffer(5230) := X"00000000";
		ram_buffer(5231) := X"28CA0008";
		ram_buffer(5232) := X"1540003E";
		ram_buffer(5233) := X"00801025";
		ram_buffer(5234) := X"10A00007";
		ram_buffer(5235) := X"00043823";
		ram_buffer(5236) := X"00000000";
		ram_buffer(5237) := X"30A500FF";
		ram_buffer(5238) := X"00055200";
		ram_buffer(5239) := X"00AA2825";
		ram_buffer(5240) := X"00055400";
		ram_buffer(5241) := X"00AA2825";
		ram_buffer(5242) := X"30EA0003";
		ram_buffer(5243) := X"11400003";
		ram_buffer(5244) := X"00CA3023";
		ram_buffer(5245) := X"A8850000";
		ram_buffer(5246) := X"008A2021";
		ram_buffer(5247) := X"30EA0004";
		ram_buffer(5248) := X"11400003";
		ram_buffer(5249) := X"00CA3023";
		ram_buffer(5250) := X"AC850000";
		ram_buffer(5251) := X"008A2021";
		ram_buffer(5252) := X"30D8003F";
		ram_buffer(5253) := X"10D80016";
		ram_buffer(5254) := X"00D83823";
		ram_buffer(5255) := X"00873821";
		ram_buffer(5256) := X"AC850000";
		ram_buffer(5257) := X"AC850004";
		ram_buffer(5258) := X"AC850008";
		ram_buffer(5259) := X"AC85000C";
		ram_buffer(5260) := X"AC850010";
		ram_buffer(5261) := X"AC850014";
		ram_buffer(5262) := X"AC850018";
		ram_buffer(5263) := X"AC85001C";
		ram_buffer(5264) := X"AC850020";
		ram_buffer(5265) := X"AC850024";
		ram_buffer(5266) := X"AC850028";
		ram_buffer(5267) := X"AC85002C";
		ram_buffer(5268) := X"AC850030";
		ram_buffer(5269) := X"AC850034";
		ram_buffer(5270) := X"AC850038";
		ram_buffer(5271) := X"AC85003C";
		ram_buffer(5272) := X"24840040";
		ram_buffer(5273) := X"1487FFEE";
		ram_buffer(5274) := X"00000000";
		ram_buffer(5275) := X"03003025";
		ram_buffer(5276) := X"30D8001F";
		ram_buffer(5277) := X"10D8000A";
		ram_buffer(5278) := X"00000000";
		ram_buffer(5279) := X"AC850000";
		ram_buffer(5280) := X"AC850004";
		ram_buffer(5281) := X"AC850008";
		ram_buffer(5282) := X"AC85000C";
		ram_buffer(5283) := X"AC850010";
		ram_buffer(5284) := X"AC850014";
		ram_buffer(5285) := X"AC850018";
		ram_buffer(5286) := X"AC85001C";
		ram_buffer(5287) := X"24840020";
		ram_buffer(5288) := X"33060003";
		ram_buffer(5289) := X"10D80005";
		ram_buffer(5290) := X"03063823";
		ram_buffer(5291) := X"00873821";
		ram_buffer(5292) := X"24840004";
		ram_buffer(5293) := X"1487FFFE";
		ram_buffer(5294) := X"AC85FFFC";
		ram_buffer(5295) := X"18C00004";
		ram_buffer(5296) := X"00863821";
		ram_buffer(5297) := X"24840001";
		ram_buffer(5298) := X"1487FFFE";
		ram_buffer(5299) := X"A085FFFF";
		ram_buffer(5300) := X"03E00008";
		ram_buffer(5301) := X"00000000";
		ram_buffer(5302) := X"24820001";
		ram_buffer(5303) := X"90830000";
		ram_buffer(5304) := X"00000000";
		ram_buffer(5305) := X"1460FFFD";
		ram_buffer(5306) := X"24840001";
		ram_buffer(5307) := X"03E00008";
		ram_buffer(5308) := X"00821023";
		ram_buffer(5309) := X"2A2A2A2A";
		ram_buffer(5310) := X"20546872";
		ram_buffer(5311) := X"6561642D";
		ram_buffer(5312) := X"4D657472";
		ram_buffer(5313) := X"69632050";
		ram_buffer(5314) := X"7265656D";
		ram_buffer(5315) := X"70746976";
		ram_buffer(5316) := X"65205363";
		ram_buffer(5317) := X"68656475";
		ram_buffer(5318) := X"6C696E67";
		ram_buffer(5319) := X"20546573";
		ram_buffer(5320) := X"74202A2A";
		ram_buffer(5321) := X"2A2A2052";
		ram_buffer(5322) := X"656C6174";
		ram_buffer(5323) := X"69766520";
		ram_buffer(5324) := X"54696D65";
		ram_buffer(5325) := X"3A202575";
		ram_buffer(5326) := X"0A0D0000";
		ram_buffer(5327) := X"4552524F";
		ram_buffer(5328) := X"523A2049";
		ram_buffer(5329) := X"6E76616C";
		ram_buffer(5330) := X"69642063";
		ram_buffer(5331) := X"6F756E74";
		ram_buffer(5332) := X"65722076";
		ram_buffer(5333) := X"616C7565";
		ram_buffer(5334) := X"2873292E";
		ram_buffer(5335) := X"20507265";
		ram_buffer(5336) := X"656D7074";
		ram_buffer(5337) := X"69766520";
		ram_buffer(5338) := X"636F756E";
		ram_buffer(5339) := X"74657273";
		ram_buffer(5340) := X"2073686F";
		ram_buffer(5341) := X"756C6420";
		ram_buffer(5342) := X"6E6F7420";
		ram_buffer(5343) := X"6265206D";
		ram_buffer(5344) := X"6F726520";
		ram_buffer(5345) := X"74686174";
		ram_buffer(5346) := X"20312064";
		ram_buffer(5347) := X"69666665";
		ram_buffer(5348) := X"72656E74";
		ram_buffer(5349) := X"20746861";
		ram_buffer(5350) := X"6E207468";
		ram_buffer(5351) := X"65206176";
		ram_buffer(5352) := X"65726167";
		ram_buffer(5353) := X"65210A0D";
		ram_buffer(5354) := X"00000000";
		ram_buffer(5355) := X"54696D65";
		ram_buffer(5356) := X"20746D5F";
		ram_buffer(5357) := X"70726565";
		ram_buffer(5358) := X"6D707469";
		ram_buffer(5359) := X"76655F74";
		ram_buffer(5360) := X"68726561";
		ram_buffer(5361) := X"645F305F";
		ram_buffer(5362) := X"636F756E";
		ram_buffer(5363) := X"74657220";
		ram_buffer(5364) := X"546F7461";
		ram_buffer(5365) := X"6C3A2020";
		ram_buffer(5366) := X"25750A0D";
		ram_buffer(5367) := X"00000000";
		ram_buffer(5368) := X"54696D65";
		ram_buffer(5369) := X"20746D5F";
		ram_buffer(5370) := X"70726565";
		ram_buffer(5371) := X"6D707469";
		ram_buffer(5372) := X"76655F74";
		ram_buffer(5373) := X"68726561";
		ram_buffer(5374) := X"645F315F";
		ram_buffer(5375) := X"636F756E";
		ram_buffer(5376) := X"74657220";
		ram_buffer(5377) := X"546F7461";
		ram_buffer(5378) := X"6C3A2020";
		ram_buffer(5379) := X"25750A0D";
		ram_buffer(5380) := X"00000000";
		ram_buffer(5381) := X"54696D65";
		ram_buffer(5382) := X"20746D5F";
		ram_buffer(5383) := X"70726565";
		ram_buffer(5384) := X"6D707469";
		ram_buffer(5385) := X"76655F74";
		ram_buffer(5386) := X"68726561";
		ram_buffer(5387) := X"645F325F";
		ram_buffer(5388) := X"636F756E";
		ram_buffer(5389) := X"74657220";
		ram_buffer(5390) := X"546F7461";
		ram_buffer(5391) := X"6C3A2020";
		ram_buffer(5392) := X"25750A0D";
		ram_buffer(5393) := X"00000000";
		ram_buffer(5394) := X"54696D65";
		ram_buffer(5395) := X"20746D5F";
		ram_buffer(5396) := X"70726565";
		ram_buffer(5397) := X"6D707469";
		ram_buffer(5398) := X"76655F74";
		ram_buffer(5399) := X"68726561";
		ram_buffer(5400) := X"645F335F";
		ram_buffer(5401) := X"636F756E";
		ram_buffer(5402) := X"74657220";
		ram_buffer(5403) := X"546F7461";
		ram_buffer(5404) := X"6C3A2020";
		ram_buffer(5405) := X"25750A0D";
		ram_buffer(5406) := X"00000000";
		ram_buffer(5407) := X"54696D65";
		ram_buffer(5408) := X"20746D5F";
		ram_buffer(5409) := X"70726565";
		ram_buffer(5410) := X"6D707469";
		ram_buffer(5411) := X"76655F74";
		ram_buffer(5412) := X"68726561";
		ram_buffer(5413) := X"645F345F";
		ram_buffer(5414) := X"636F756E";
		ram_buffer(5415) := X"74657220";
		ram_buffer(5416) := X"546F7461";
		ram_buffer(5417) := X"6C3A2020";
		ram_buffer(5418) := X"25750A0D";
		ram_buffer(5419) := X"00000000";
		ram_buffer(5420) := X"54696D65";
		ram_buffer(5421) := X"20506572";
		ram_buffer(5422) := X"696F6420";
		ram_buffer(5423) := X"546F7461";
		ram_buffer(5424) := X"6C3A2020";
		ram_buffer(5425) := X"25750A0D";
		ram_buffer(5426) := X"0A0D0000";
		ram_buffer(5427) := X"416C6976";
		ram_buffer(5428) := X"652E2E2E";
		ram_buffer(5429) := X"0A0D0000";
		ram_buffer(5430) := X"41737365";
		ram_buffer(5431) := X"72743A0A";
		ram_buffer(5432) := X"0D4D6573";
		ram_buffer(5433) := X"73616765";
		ram_buffer(5434) := X"3A25730A";
		ram_buffer(5435) := X"0D4C696E";
		ram_buffer(5436) := X"653A2564";
		ram_buffer(5437) := X"0A0D0000";
		ram_buffer(5438) := X"746D5F70";
		ram_buffer(5439) := X"6F727469";
		ram_buffer(5440) := X"6E675F6C";
		ram_buffer(5441) := X"61796572";
		ram_buffer(5442) := X"5F667265";
		ram_buffer(5443) := X"6572746F";
		ram_buffer(5444) := X"732E6300";
		ram_buffer(5445) := X"2E2E2F2E";
		ram_buffer(5446) := X"2E2F6672";
		ram_buffer(5447) := X"65657274";
		ram_buffer(5448) := X"6F732F71";
		ram_buffer(5449) := X"75657565";
		ram_buffer(5450) := X"2E630000";
		ram_buffer(5451) := X"2E2E2F2E";
		ram_buffer(5452) := X"2E2F6672";
		ram_buffer(5453) := X"65657274";
		ram_buffer(5454) := X"6F732F74";
		ram_buffer(5455) := X"61736B73";
		ram_buffer(5456) := X"2E630000";
		ram_buffer(5457) := X"49444C45";
		ram_buffer(5458) := X"00000000";
		ram_buffer(5459) := X"2E2E2F2E";
		ram_buffer(5460) := X"2E2F6672";
		ram_buffer(5461) := X"65657274";
		ram_buffer(5462) := X"6F732F70";
		ram_buffer(5463) := X"6F72742E";
		ram_buffer(5464) := X"63000000";
		ram_buffer(5465) := X"2E2E2F2E";
		ram_buffer(5466) := X"2E2F6672";
		ram_buffer(5467) := X"65657274";
		ram_buffer(5468) := X"6F732F68";
		ram_buffer(5469) := X"6561705F";
		ram_buffer(5470) := X"342E6300";
		ram_buffer(5471) := X"00000000";
		ram_buffer(5472) := X"00000100";
		ram_buffer(5473) := X"01010001";
		ram_buffer(5474) := X"00000000";
		ram_buffer(5475) := X"00000000";
		ram_buffer(5476) := X"00000000";
		ram_buffer(5477) := X"00000000";
		return ram_buffer;
	end;
end;
