library ieee;
use ieee.std_logic_1164.all;

package bram_pack is

	constant cpu_width : integer := 32;
	constant ram_size : integer := 16384;
	subtype word_type is std_logic_vector(cpu_width-1 downto 0);
	type ram_type is array(0 to ram_size-1) of word_type;
	function load_hex return ram_type;

end package;

package body bram_pack is

	function load_hex return ram_type is
		variable ram_buffer : ram_type := (others=>(others=>'0'));
	begin
		ram_buffer(0) := X"3C1C0001";
		ram_buffer(1) := X"279C83F0";
		ram_buffer(2) := X"3C050000";
		ram_buffer(3) := X"24A503FC";
		ram_buffer(4) := X"3C040000";
		ram_buffer(5) := X"24840654";
		ram_buffer(6) := X"3C1D0000";
		ram_buffer(7) := X"27BD05F8";
		ram_buffer(8) := X"ACA00000";
		ram_buffer(9) := X"00A4182A";
		ram_buffer(10) := X"1460FFFD";
		ram_buffer(11) := X"24A50004";
		ram_buffer(12) := X"0C00007C";
		ram_buffer(13) := X"00000000";
		ram_buffer(14) := X"0800000E";
		ram_buffer(15) := X"23BDFF98";
		ram_buffer(16) := X"AFA10010";
		ram_buffer(17) := X"AFA20014";
		ram_buffer(18) := X"AFA30018";
		ram_buffer(19) := X"AFA4001C";
		ram_buffer(20) := X"AFA50020";
		ram_buffer(21) := X"AFA60024";
		ram_buffer(22) := X"AFA70028";
		ram_buffer(23) := X"AFA8002C";
		ram_buffer(24) := X"AFA90030";
		ram_buffer(25) := X"AFAA0034";
		ram_buffer(26) := X"AFAB0038";
		ram_buffer(27) := X"AFAC003C";
		ram_buffer(28) := X"AFAD0040";
		ram_buffer(29) := X"AFAE0044";
		ram_buffer(30) := X"AFAF0048";
		ram_buffer(31) := X"AFB8004C";
		ram_buffer(32) := X"AFB90050";
		ram_buffer(33) := X"AFBF0054";
		ram_buffer(34) := X"401A7000";
		ram_buffer(35) := X"235AFFFC";
		ram_buffer(36) := X"AFBA0058";
		ram_buffer(37) := X"0000D810";
		ram_buffer(38) := X"AFBB005C";
		ram_buffer(39) := X"0000D812";
		ram_buffer(40) := X"AFBB0060";
		ram_buffer(41) := X"0C0000CC";
		ram_buffer(42) := X"23A50000";
		ram_buffer(43) := X"8FA10010";
		ram_buffer(44) := X"8FA20014";
		ram_buffer(45) := X"8FA30018";
		ram_buffer(46) := X"8FA4001C";
		ram_buffer(47) := X"8FA50020";
		ram_buffer(48) := X"8FA60024";
		ram_buffer(49) := X"8FA70028";
		ram_buffer(50) := X"8FA8002C";
		ram_buffer(51) := X"8FA90030";
		ram_buffer(52) := X"8FAA0034";
		ram_buffer(53) := X"8FAB0038";
		ram_buffer(54) := X"8FAC003C";
		ram_buffer(55) := X"8FAD0040";
		ram_buffer(56) := X"8FAE0044";
		ram_buffer(57) := X"8FAF0048";
		ram_buffer(58) := X"8FB8004C";
		ram_buffer(59) := X"8FB90050";
		ram_buffer(60) := X"8FBF0054";
		ram_buffer(61) := X"8FBA0058";
		ram_buffer(62) := X"8FBB005C";
		ram_buffer(63) := X"03600011";
		ram_buffer(64) := X"8FBB0060";
		ram_buffer(65) := X"03600013";
		ram_buffer(66) := X"23BD0068";
		ram_buffer(67) := X"341B0001";
		ram_buffer(68) := X"03400008";
		ram_buffer(69) := X"409B6000";
		ram_buffer(70) := X"40026000";
		ram_buffer(71) := X"03E00008";
		ram_buffer(72) := X"40846000";
		ram_buffer(73) := X"3C050000";
		ram_buffer(74) := X"24A50150";
		ram_buffer(75) := X"8CA60000";
		ram_buffer(76) := X"AC06003C";
		ram_buffer(77) := X"8CA60004";
		ram_buffer(78) := X"AC060040";
		ram_buffer(79) := X"8CA60008";
		ram_buffer(80) := X"AC060044";
		ram_buffer(81) := X"8CA6000C";
		ram_buffer(82) := X"03E00008";
		ram_buffer(83) := X"AC060048";
		ram_buffer(84) := X"3C1A1000";
		ram_buffer(85) := X"375A003C";
		ram_buffer(86) := X"03400008";
		ram_buffer(87) := X"00000000";
		ram_buffer(88) := X"AC900000";
		ram_buffer(89) := X"AC910004";
		ram_buffer(90) := X"AC920008";
		ram_buffer(91) := X"AC93000C";
		ram_buffer(92) := X"AC940010";
		ram_buffer(93) := X"AC950014";
		ram_buffer(94) := X"AC960018";
		ram_buffer(95) := X"AC97001C";
		ram_buffer(96) := X"AC9E0020";
		ram_buffer(97) := X"AC9C0024";
		ram_buffer(98) := X"AC9D0028";
		ram_buffer(99) := X"AC9F002C";
		ram_buffer(100) := X"03E00008";
		ram_buffer(101) := X"34020000";
		ram_buffer(102) := X"8C900000";
		ram_buffer(103) := X"8C910004";
		ram_buffer(104) := X"8C920008";
		ram_buffer(105) := X"8C93000C";
		ram_buffer(106) := X"8C940010";
		ram_buffer(107) := X"8C950014";
		ram_buffer(108) := X"8C960018";
		ram_buffer(109) := X"8C97001C";
		ram_buffer(110) := X"8C9E0020";
		ram_buffer(111) := X"8C9C0024";
		ram_buffer(112) := X"8C9D0028";
		ram_buffer(113) := X"8C9F002C";
		ram_buffer(114) := X"03E00008";
		ram_buffer(115) := X"34A20000";
		ram_buffer(116) := X"00850019";
		ram_buffer(117) := X"00001012";
		ram_buffer(118) := X"00002010";
		ram_buffer(119) := X"03E00008";
		ram_buffer(120) := X"ACC40000";
		ram_buffer(121) := X"0000000C";
		ram_buffer(122) := X"03E00008";
		ram_buffer(123) := X"00000000";
		ram_buffer(124) := X"27BDFFE8";
		ram_buffer(125) := X"3C0344A0";
		ram_buffer(126) := X"AFB00010";
		ram_buffer(127) := X"3C100000";
		ram_buffer(128) := X"AE030610";
		ram_buffer(129) := X"3C0344A2";
		ram_buffer(130) := X"AF838014";
		ram_buffer(131) := X"3C03017D";
		ram_buffer(132) := X"3C0444A1";
		ram_buffer(133) := X"24637840";
		ram_buffer(134) := X"AFBF0014";
		ram_buffer(135) := X"AF848010";
		ram_buffer(136) := X"AC830004";
		ram_buffer(137) := X"3C030000";
		ram_buffer(138) := X"26020610";
		ram_buffer(139) := X"24630304";
		ram_buffer(140) := X"AC43000C";
		ram_buffer(141) := X"3C030000";
		ram_buffer(142) := X"246302DC";
		ram_buffer(143) := X"24040001";
		ram_buffer(144) := X"AC430004";
		ram_buffer(145) := X"AC400014";
		ram_buffer(146) := X"AC40001C";
		ram_buffer(147) := X"AC400024";
		ram_buffer(148) := X"AC40002C";
		ram_buffer(149) := X"AC400034";
		ram_buffer(150) := X"AC40003C";
		ram_buffer(151) := X"AC400010";
		ram_buffer(152) := X"0C000046";
		ram_buffer(153) := X"AC400008";
		ram_buffer(154) := X"8E020610";
		ram_buffer(155) := X"240300FF";
		ram_buffer(156) := X"AC430000";
		ram_buffer(157) := X"8F828010";
		ram_buffer(158) := X"24030003";
		ram_buffer(159) := X"AC430000";
		ram_buffer(160) := X"8F828014";
		ram_buffer(161) := X"24030001";
		ram_buffer(162) := X"AC430000";
		ram_buffer(163) := X"240400FF";
		ram_buffer(164) := X"8F828008";
		ram_buffer(165) := X"00000000";
		ram_buffer(166) := X"1040FFFD";
		ram_buffer(167) := X"00000000";
		ram_buffer(168) := X"8E020610";
		ram_buffer(169) := X"00000000";
		ram_buffer(170) := X"AC400000";
		ram_buffer(171) := X"AF808008";
		ram_buffer(172) := X"8F828018";
		ram_buffer(173) := X"8F83800C";
		ram_buffer(174) := X"00000000";
		ram_buffer(175) := X"00430018";
		ram_buffer(176) := X"8F838014";
		ram_buffer(177) := X"00001012";
		ram_buffer(178) := X"AC620008";
		ram_buffer(179) := X"8E020610";
		ram_buffer(180) := X"00000000";
		ram_buffer(181) := X"1000FFEE";
		ram_buffer(182) := X"AC440000";
		ram_buffer(183) := X"8F82800C";
		ram_buffer(184) := X"00000000";
		ram_buffer(185) := X"2C420001";
		ram_buffer(186) := X"AF82800C";
		ram_buffer(187) := X"24020001";
		ram_buffer(188) := X"AF828008";
		ram_buffer(189) := X"8F828010";
		ram_buffer(190) := X"24030007";
		ram_buffer(191) := X"03E00008";
		ram_buffer(192) := X"AC430000";
		ram_buffer(193) := X"8F838014";
		ram_buffer(194) := X"24020001";
		ram_buffer(195) := X"8C630004";
		ram_buffer(196) := X"00000000";
		ram_buffer(197) := X"AF838018";
		ram_buffer(198) := X"AF82800C";
		ram_buffer(199) := X"AF828008";
		ram_buffer(200) := X"8F828014";
		ram_buffer(201) := X"24030003";
		ram_buffer(202) := X"03E00008";
		ram_buffer(203) := X"AC430000";
		ram_buffer(204) := X"27BDFFE0";
		ram_buffer(205) := X"AFB10018";
		ram_buffer(206) := X"3C110000";
		ram_buffer(207) := X"8E220610";
		ram_buffer(208) := X"AFBF001C";
		ram_buffer(209) := X"8C420004";
		ram_buffer(210) := X"00000000";
		ram_buffer(211) := X"2C430008";
		ram_buffer(212) := X"10600010";
		ram_buffer(213) := X"AFB00014";
		ram_buffer(214) := X"3C100000";
		ram_buffer(215) := X"26100614";
		ram_buffer(216) := X"000210C0";
		ram_buffer(217) := X"02021021";
		ram_buffer(218) := X"8C430000";
		ram_buffer(219) := X"8C440004";
		ram_buffer(220) := X"0060F809";
		ram_buffer(221) := X"00000000";
		ram_buffer(222) := X"8E220610";
		ram_buffer(223) := X"00000000";
		ram_buffer(224) := X"8C420004";
		ram_buffer(225) := X"00000000";
		ram_buffer(226) := X"2C430008";
		ram_buffer(227) := X"1460FFF4";
		ram_buffer(228) := X"00000000";
		ram_buffer(229) := X"8FBF001C";
		ram_buffer(230) := X"8FB10018";
		ram_buffer(231) := X"8FB00014";
		ram_buffer(232) := X"03E00008";
		ram_buffer(233) := X"27BD0020";
		ram_buffer(234) := X"10C00011";
		ram_buffer(235) := X"00C51821";
		ram_buffer(236) := X"2406FFE0";
		ram_buffer(237) := X"00661024";
		ram_buffer(238) := X"0043182B";
		ram_buffer(239) := X"00031940";
		ram_buffer(240) := X"24420020";
		ram_buffer(241) := X"00A62824";
		ram_buffer(242) := X"00431821";
		ram_buffer(243) := X"10A30008";
		ram_buffer(244) := X"3C021000";
		ram_buffer(245) := X"00822021";
		ram_buffer(246) := X"00A61024";
		ram_buffer(247) := X"AC820000";
		ram_buffer(248) := X"AC400000";
		ram_buffer(249) := X"24A50020";
		ram_buffer(250) := X"14A3FFFC";
		ram_buffer(251) := X"00A61024";
		ram_buffer(252) := X"03E00008";
		ram_buffer(253) := X"00000000";
		ram_buffer(254) := X"00000001";
		ram_buffer(255) := X"00000000";
		ram_buffer(256) := X"00000000";
		ram_buffer(257) := X"00000000";
		ram_buffer(258) := X"00000000";
		ram_buffer(259) := X"00000000";
		ram_buffer(260) := X"00000000";
		ram_buffer(261) := X"00000000";
		ram_buffer(262) := X"00000000";
		ram_buffer(263) := X"00000000";
		ram_buffer(264) := X"00000000";
		ram_buffer(265) := X"00000000";
		ram_buffer(266) := X"00000000";
		ram_buffer(267) := X"00000000";
		ram_buffer(268) := X"00000000";
		ram_buffer(269) := X"00000000";
		ram_buffer(270) := X"00000000";
		ram_buffer(271) := X"00000000";
		ram_buffer(272) := X"00000000";
		ram_buffer(273) := X"00000000";
		ram_buffer(274) := X"00000000";

		return ram_buffer;
	end;
end;
