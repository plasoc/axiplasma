----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 01/28/2017 04:46:42 PM
-- Design Name: 
-- Module Name: plasoc_int_axi4_read_cntrl - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use work.mlitesoc_pack.all;

entity plasoc_int_axi4_read_cntrl is
--  Port ( );
end plasoc_int_axi4_read_cntrl;

architecture Behavioral of plasoc_int_axi4_read_cntrl is

begin


end Behavioral;
