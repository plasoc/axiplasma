
library ieee;
use ieee.std_logic_1164.all;

package vc707_pack is

    constant vc707_default_gpio_width : integer := 8;
    
end package;

