library ieee;
use ieee.std_logic_1164.all;

package bram_pack is

	constant cpu_width : integer := 32;
	constant ram_size : integer := 8192;
	subtype word_type is std_logic_vector(cpu_width-1 downto 0);
	type ram_type is array(0 to ram_size-1) of word_type;
	function load_hex return ram_type;

end package;

package body bram_pack is

	function load_hex return ram_type is
		variable ram_buffer : ram_type := (others=>(others=>'0'));
	begin
		ram_buffer(0) := X"3C1C0001";
		ram_buffer(1) := X"279CC610";
		ram_buffer(2) := X"3C050000";
		ram_buffer(3) := X"24A5461C";
		ram_buffer(4) := X"3C040000";
		ram_buffer(5) := X"24846A24";
		ram_buffer(6) := X"3C1D0000";
		ram_buffer(7) := X"27BD6938";
		ram_buffer(8) := X"ACA00000";
		ram_buffer(9) := X"00A4182A";
		ram_buffer(10) := X"1460FFFD";
		ram_buffer(11) := X"24A50004";
		ram_buffer(12) := X"0C00007C";
		ram_buffer(13) := X"00000000";
		ram_buffer(14) := X"0800000E";
		ram_buffer(15) := X"23BDFF98";
		ram_buffer(16) := X"AFA10010";
		ram_buffer(17) := X"AFA20014";
		ram_buffer(18) := X"AFA30018";
		ram_buffer(19) := X"AFA4001C";
		ram_buffer(20) := X"AFA50020";
		ram_buffer(21) := X"AFA60024";
		ram_buffer(22) := X"AFA70028";
		ram_buffer(23) := X"AFA8002C";
		ram_buffer(24) := X"AFA90030";
		ram_buffer(25) := X"AFAA0034";
		ram_buffer(26) := X"AFAB0038";
		ram_buffer(27) := X"AFAC003C";
		ram_buffer(28) := X"AFAD0040";
		ram_buffer(29) := X"AFAE0044";
		ram_buffer(30) := X"AFAF0048";
		ram_buffer(31) := X"AFB8004C";
		ram_buffer(32) := X"AFB90050";
		ram_buffer(33) := X"AFBF0054";
		ram_buffer(34) := X"401A7000";
		ram_buffer(35) := X"235AFFFC";
		ram_buffer(36) := X"AFBA0058";
		ram_buffer(37) := X"0000D810";
		ram_buffer(38) := X"AFBB005C";
		ram_buffer(39) := X"0000D812";
		ram_buffer(40) := X"AFBB0060";
		ram_buffer(41) := X"0C000FF6";
		ram_buffer(42) := X"23A50000";
		ram_buffer(43) := X"8FA10010";
		ram_buffer(44) := X"8FA20014";
		ram_buffer(45) := X"8FA30018";
		ram_buffer(46) := X"8FA4001C";
		ram_buffer(47) := X"8FA50020";
		ram_buffer(48) := X"8FA60024";
		ram_buffer(49) := X"8FA70028";
		ram_buffer(50) := X"8FA8002C";
		ram_buffer(51) := X"8FA90030";
		ram_buffer(52) := X"8FAA0034";
		ram_buffer(53) := X"8FAB0038";
		ram_buffer(54) := X"8FAC003C";
		ram_buffer(55) := X"8FAD0040";
		ram_buffer(56) := X"8FAE0044";
		ram_buffer(57) := X"8FAF0048";
		ram_buffer(58) := X"8FB8004C";
		ram_buffer(59) := X"8FB90050";
		ram_buffer(60) := X"8FBF0054";
		ram_buffer(61) := X"8FBA0058";
		ram_buffer(62) := X"8FBB005C";
		ram_buffer(63) := X"03600011";
		ram_buffer(64) := X"8FBB0060";
		ram_buffer(65) := X"03600013";
		ram_buffer(66) := X"23BD0068";
		ram_buffer(67) := X"341B0001";
		ram_buffer(68) := X"03400008";
		ram_buffer(69) := X"409B6000";
		ram_buffer(70) := X"40026000";
		ram_buffer(71) := X"03E00008";
		ram_buffer(72) := X"40846000";
		ram_buffer(73) := X"3C050000";
		ram_buffer(74) := X"24A50150";
		ram_buffer(75) := X"8CA60000";
		ram_buffer(76) := X"AC06003C";
		ram_buffer(77) := X"8CA60004";
		ram_buffer(78) := X"AC060040";
		ram_buffer(79) := X"8CA60008";
		ram_buffer(80) := X"AC060044";
		ram_buffer(81) := X"8CA6000C";
		ram_buffer(82) := X"03E00008";
		ram_buffer(83) := X"AC060048";
		ram_buffer(84) := X"3C1A1000";
		ram_buffer(85) := X"375A003C";
		ram_buffer(86) := X"03400008";
		ram_buffer(87) := X"00000000";
		ram_buffer(88) := X"AC900000";
		ram_buffer(89) := X"AC910004";
		ram_buffer(90) := X"AC920008";
		ram_buffer(91) := X"AC93000C";
		ram_buffer(92) := X"AC940010";
		ram_buffer(93) := X"AC950014";
		ram_buffer(94) := X"AC960018";
		ram_buffer(95) := X"AC97001C";
		ram_buffer(96) := X"AC9E0020";
		ram_buffer(97) := X"AC9C0024";
		ram_buffer(98) := X"AC9D0028";
		ram_buffer(99) := X"AC9F002C";
		ram_buffer(100) := X"03E00008";
		ram_buffer(101) := X"34020000";
		ram_buffer(102) := X"8C900000";
		ram_buffer(103) := X"8C910004";
		ram_buffer(104) := X"8C920008";
		ram_buffer(105) := X"8C93000C";
		ram_buffer(106) := X"8C940010";
		ram_buffer(107) := X"8C950014";
		ram_buffer(108) := X"8C960018";
		ram_buffer(109) := X"8C97001C";
		ram_buffer(110) := X"8C9E0020";
		ram_buffer(111) := X"8C9C0024";
		ram_buffer(112) := X"8C9D0028";
		ram_buffer(113) := X"8C9F002C";
		ram_buffer(114) := X"03E00008";
		ram_buffer(115) := X"34A20000";
		ram_buffer(116) := X"00850019";
		ram_buffer(117) := X"00001012";
		ram_buffer(118) := X"00002010";
		ram_buffer(119) := X"03E00008";
		ram_buffer(120) := X"ACC40000";
		ram_buffer(121) := X"0000000C";
		ram_buffer(122) := X"03E00008";
		ram_buffer(123) := X"00000000";
		ram_buffer(124) := X"27BDFFD0";
		ram_buffer(125) := X"00002025";
		ram_buffer(126) := X"AFB0001C";
		ram_buffer(127) := X"AFBF002C";
		ram_buffer(128) := X"AFB30028";
		ram_buffer(129) := X"AFB20024";
		ram_buffer(130) := X"AFB10020";
		ram_buffer(131) := X"0C000046";
		ram_buffer(132) := X"3C100000";
		ram_buffer(133) := X"3C0244A0";
		ram_buffer(134) := X"AE026950";
		ram_buffer(135) := X"3C030000";
		ram_buffer(136) := X"3C020000";
		ram_buffer(137) := X"24426954";
		ram_buffer(138) := X"24636994";
		ram_buffer(139) := X"24420008";
		ram_buffer(140) := X"1443FFFE";
		ram_buffer(141) := X"AC40FFF8";
		ram_buffer(142) := X"3C0244A2";
		ram_buffer(143) := X"3C030000";
		ram_buffer(144) := X"AF82805C";
		ram_buffer(145) := X"24630654";
		ram_buffer(146) := X"26026950";
		ram_buffer(147) := X"AC43000C";
		ram_buffer(148) := X"3404C350";
		ram_buffer(149) := X"3C0344A1";
		ram_buffer(150) := X"AF838058";
		ram_buffer(151) := X"AC400010";
		ram_buffer(152) := X"AC640004";
		ram_buffer(153) := X"3C030000";
		ram_buffer(154) := X"24630620";
		ram_buffer(155) := X"3C040000";
		ram_buffer(156) := X"AC430004";
		ram_buffer(157) := X"24060040";
		ram_buffer(158) := X"00002825";
		ram_buffer(159) := X"24846994";
		ram_buffer(160) := X"0C001119";
		ram_buffer(161) := X"AC400008";
		ram_buffer(162) := X"00003025";
		ram_buffer(163) := X"24050004";
		ram_buffer(164) := X"0C000361";
		ram_buffer(165) := X"24040008";
		ram_buffer(166) := X"14400006";
		ram_buffer(167) := X"AF828064";
		ram_buffer(168) := X"8F82805C";
		ram_buffer(169) := X"240300B2";
		ram_buffer(170) := X"AC430008";
		ram_buffer(171) := X"1000FFFF";
		ram_buffer(172) := X"00000000";
		ram_buffer(173) := X"00002825";
		ram_buffer(174) := X"0C000385";
		ram_buffer(175) := X"24040008";
		ram_buffer(176) := X"14400006";
		ram_buffer(177) := X"AF828060";
		ram_buffer(178) := X"8F82805C";
		ram_buffer(179) := X"240300B4";
		ram_buffer(180) := X"AC430008";
		ram_buffer(181) := X"1000FFFF";
		ram_buffer(182) := X"00000000";
		ram_buffer(183) := X"24110003";
		ram_buffer(184) := X"3C050000";
		ram_buffer(185) := X"3C040000";
		ram_buffer(186) := X"AFA00014";
		ram_buffer(187) := X"AFB10010";
		ram_buffer(188) := X"00003825";
		ram_buffer(189) := X"2406012C";
		ram_buffer(190) := X"24A5459C";
		ram_buffer(191) := X"0C000A44";
		ram_buffer(192) := X"24840714";
		ram_buffer(193) := X"00409825";
		ram_buffer(194) := X"24020001";
		ram_buffer(195) := X"12620006";
		ram_buffer(196) := X"240300B6";
		ram_buffer(197) := X"8F82805C";
		ram_buffer(198) := X"00000000";
		ram_buffer(199) := X"AC430008";
		ram_buffer(200) := X"1000FFFF";
		ram_buffer(201) := X"00000000";
		ram_buffer(202) := X"27828068";
		ram_buffer(203) := X"3C050000";
		ram_buffer(204) := X"3C040000";
		ram_buffer(205) := X"AFA20014";
		ram_buffer(206) := X"AFB10010";
		ram_buffer(207) := X"00003825";
		ram_buffer(208) := X"2406012C";
		ram_buffer(209) := X"24A545A4";
		ram_buffer(210) := X"0C000A44";
		ram_buffer(211) := X"2484069C";
		ram_buffer(212) := X"10530006";
		ram_buffer(213) := X"00409025";
		ram_buffer(214) := X"8F82805C";
		ram_buffer(215) := X"240300B8";
		ram_buffer(216) := X"AC430008";
		ram_buffer(217) := X"1000FFFF";
		ram_buffer(218) := X"00000000";
		ram_buffer(219) := X"3C050000";
		ram_buffer(220) := X"3C040000";
		ram_buffer(221) := X"AFA00014";
		ram_buffer(222) := X"AFB10010";
		ram_buffer(223) := X"00003825";
		ram_buffer(224) := X"2406012C";
		ram_buffer(225) := X"24A545AC";
		ram_buffer(226) := X"0C000A44";
		ram_buffer(227) := X"248406D8";
		ram_buffer(228) := X"10520006";
		ram_buffer(229) := X"240300BA";
		ram_buffer(230) := X"8F82805C";
		ram_buffer(231) := X"00000000";
		ram_buffer(232) := X"AC430008";
		ram_buffer(233) := X"1000FFFF";
		ram_buffer(234) := X"00000000";
		ram_buffer(235) := X"8E036950";
		ram_buffer(236) := X"240400FF";
		ram_buffer(237) := X"AC640000";
		ram_buffer(238) := X"8F838058";
		ram_buffer(239) := X"00000000";
		ram_buffer(240) := X"AC710000";
		ram_buffer(241) := X"8F83805C";
		ram_buffer(242) := X"00000000";
		ram_buffer(243) := X"0C000AFF";
		ram_buffer(244) := X"AC620000";
		ram_buffer(245) := X"8F82805C";
		ram_buffer(246) := X"240300C6";
		ram_buffer(247) := X"AC430008";
		ram_buffer(248) := X"1000FFFF";
		ram_buffer(249) := X"00000000";
		ram_buffer(250) := X"2082FF98";
		ram_buffer(251) := X"AC450058";
		ram_buffer(252) := X"03E00008";
		ram_buffer(253) := X"AC46001C";
		ram_buffer(254) := X"3C1A0000";
		ram_buffer(255) := X"375A4664";
		ram_buffer(256) := X"8F5B0000";
		ram_buffer(257) := X"AF400000";
		ram_buffer(258) := X"23BDFF98";
		ram_buffer(259) := X"AFA10010";
		ram_buffer(260) := X"AFA20014";
		ram_buffer(261) := X"AFA30018";
		ram_buffer(262) := X"AFA4001C";
		ram_buffer(263) := X"AFA50020";
		ram_buffer(264) := X"AFA60024";
		ram_buffer(265) := X"AFA70028";
		ram_buffer(266) := X"AFA8002C";
		ram_buffer(267) := X"AFA90030";
		ram_buffer(268) := X"AFAA0034";
		ram_buffer(269) := X"AFAB0038";
		ram_buffer(270) := X"AFAC003C";
		ram_buffer(271) := X"AFAD0040";
		ram_buffer(272) := X"AFAE0044";
		ram_buffer(273) := X"AFAF0048";
		ram_buffer(274) := X"AFB8004C";
		ram_buffer(275) := X"AFB90050";
		ram_buffer(276) := X"AFBF0054";
		ram_buffer(277) := X"401A7000";
		ram_buffer(278) := X"17600003";
		ram_buffer(279) := X"235AFFFC";
		ram_buffer(280) := X"0800011B";
		ram_buffer(281) := X"00000000";
		ram_buffer(282) := X"235A0004";
		ram_buffer(283) := X"AFBA0058";
		ram_buffer(284) := X"0000D810";
		ram_buffer(285) := X"AFBB005C";
		ram_buffer(286) := X"0000D812";
		ram_buffer(287) := X"AFBB0060";
		ram_buffer(288) := X"3C1A0000";
		ram_buffer(289) := X"375A461C";
		ram_buffer(290) := X"8F5A0000";
		ram_buffer(291) := X"AF5D0000";
		ram_buffer(292) := X"3C1A0000";
		ram_buffer(293) := X"375A6750";
		ram_buffer(294) := X"8F5D0000";
		ram_buffer(295) := X"0C00020C";
		ram_buffer(296) := X"00000000";
		ram_buffer(297) := X"3C1A0000";
		ram_buffer(298) := X"375A6750";
		ram_buffer(299) := X"AF5D0000";
		ram_buffer(300) := X"3C1A0000";
		ram_buffer(301) := X"375A461C";
		ram_buffer(302) := X"8F5A0000";
		ram_buffer(303) := X"8F5D0000";
		ram_buffer(304) := X"8FA10010";
		ram_buffer(305) := X"8FA20014";
		ram_buffer(306) := X"8FA30018";
		ram_buffer(307) := X"8FA4001C";
		ram_buffer(308) := X"8FA50020";
		ram_buffer(309) := X"8FA60024";
		ram_buffer(310) := X"8FA70028";
		ram_buffer(311) := X"8FA8002C";
		ram_buffer(312) := X"8FA90030";
		ram_buffer(313) := X"8FAA0034";
		ram_buffer(314) := X"8FAB0038";
		ram_buffer(315) := X"8FAC003C";
		ram_buffer(316) := X"8FAD0040";
		ram_buffer(317) := X"8FAE0044";
		ram_buffer(318) := X"8FAF0048";
		ram_buffer(319) := X"8FB8004C";
		ram_buffer(320) := X"8FB90050";
		ram_buffer(321) := X"8FBF0054";
		ram_buffer(322) := X"8FBA0058";
		ram_buffer(323) := X"8FBB005C";
		ram_buffer(324) := X"03600011";
		ram_buffer(325) := X"8FBB0060";
		ram_buffer(326) := X"03600013";
		ram_buffer(327) := X"23BD0068";
		ram_buffer(328) := X"341B0001";
		ram_buffer(329) := X"03400008";
		ram_buffer(330) := X"409B6000";
		ram_buffer(331) := X"00000000";
		ram_buffer(332) := X"3C080000";
		ram_buffer(333) := X"2508055C";
		ram_buffer(334) := X"8D090000";
		ram_buffer(335) := X"AC09003C";
		ram_buffer(336) := X"8D090004";
		ram_buffer(337) := X"AC090040";
		ram_buffer(338) := X"8D090008";
		ram_buffer(339) := X"AC090044";
		ram_buffer(340) := X"8D09000C";
		ram_buffer(341) := X"03E00008";
		ram_buffer(342) := X"AC090048";
		ram_buffer(343) := X"3C1A0000";
		ram_buffer(344) := X"375A03F8";
		ram_buffer(345) := X"03400008";
		ram_buffer(346) := X"00000000";
		ram_buffer(347) := X"3C1A0000";
		ram_buffer(348) := X"375A6750";
		ram_buffer(349) := X"AF5D0000";
		ram_buffer(350) := X"3C1A0000";
		ram_buffer(351) := X"375A461C";
		ram_buffer(352) := X"8F5A0000";
		ram_buffer(353) := X"8F5D0000";
		ram_buffer(354) := X"8FA10010";
		ram_buffer(355) := X"8FA20014";
		ram_buffer(356) := X"8FA30018";
		ram_buffer(357) := X"8FA4001C";
		ram_buffer(358) := X"8FA50020";
		ram_buffer(359) := X"8FA60024";
		ram_buffer(360) := X"8FA70028";
		ram_buffer(361) := X"8FA8002C";
		ram_buffer(362) := X"8FA90030";
		ram_buffer(363) := X"8FAA0034";
		ram_buffer(364) := X"8FAB0038";
		ram_buffer(365) := X"8FAC003C";
		ram_buffer(366) := X"8FAD0040";
		ram_buffer(367) := X"8FAE0044";
		ram_buffer(368) := X"8FAF0048";
		ram_buffer(369) := X"8FB8004C";
		ram_buffer(370) := X"8FB90050";
		ram_buffer(371) := X"8FBF0054";
		ram_buffer(372) := X"8FBA0058";
		ram_buffer(373) := X"8FBB005C";
		ram_buffer(374) := X"03600011";
		ram_buffer(375) := X"8FBB0060";
		ram_buffer(376) := X"03600013";
		ram_buffer(377) := X"23BD0068";
		ram_buffer(378) := X"341B0001";
		ram_buffer(379) := X"03400008";
		ram_buffer(380) := X"409B6000";
		ram_buffer(381) := X"40806000";
		ram_buffer(382) := X"20090001";
		ram_buffer(383) := X"3C080000";
		ram_buffer(384) := X"35084664";
		ram_buffer(385) := X"AD090000";
		ram_buffer(386) := X"3C080000";
		ram_buffer(387) := X"35084658";
		ram_buffer(388) := X"AD090000";
		ram_buffer(389) := X"0000000C";
		ram_buffer(390) := X"03E00008";
		ram_buffer(391) := X"00000000";
		ram_buffer(392) := X"27BDFFE8";
		ram_buffer(393) := X"AFBF0014";
		ram_buffer(394) := X"0C000808";
		ram_buffer(395) := X"00000000";
		ram_buffer(396) := X"10400002";
		ram_buffer(397) := X"24020001";
		ram_buffer(398) := X"AF828048";
		ram_buffer(399) := X"8FBF0014";
		ram_buffer(400) := X"8F828058";
		ram_buffer(401) := X"24030007";
		ram_buffer(402) := X"AC430000";
		ram_buffer(403) := X"03E00008";
		ram_buffer(404) := X"27BD0018";
		ram_buffer(405) := X"27BDFFE0";
		ram_buffer(406) := X"AFBF001C";
		ram_buffer(407) := X"AFA00010";
		ram_buffer(408) := X"8F82805C";
		ram_buffer(409) := X"24030003";
		ram_buffer(410) := X"8F848068";
		ram_buffer(411) := X"AC430000";
		ram_buffer(412) := X"0C000F94";
		ram_buffer(413) := X"27A50010";
		ram_buffer(414) := X"8FA20010";
		ram_buffer(415) := X"00000000";
		ram_buffer(416) := X"10400002";
		ram_buffer(417) := X"24020001";
		ram_buffer(418) := X"AF828048";
		ram_buffer(419) := X"8FBF001C";
		ram_buffer(420) := X"00000000";
		ram_buffer(421) := X"03E00008";
		ram_buffer(422) := X"27BD0020";
		ram_buffer(423) := X"27BDFFE0";
		ram_buffer(424) := X"AFBF001C";
		ram_buffer(425) := X"2405FFFF";
		ram_buffer(426) := X"0C000E42";
		ram_buffer(427) := X"24040001";
		ram_buffer(428) := X"8F82805C";
		ram_buffer(429) := X"8F848064";
		ram_buffer(430) := X"8C420004";
		ram_buffer(431) := X"00003825";
		ram_buffer(432) := X"2406FFFF";
		ram_buffer(433) := X"27A50010";
		ram_buffer(434) := X"0C0003A3";
		ram_buffer(435) := X"AFA20010";
		ram_buffer(436) := X"1000FFF5";
		ram_buffer(437) := X"2405FFFF";
		ram_buffer(438) := X"27BDFFE0";
		ram_buffer(439) := X"AFBF001C";
		ram_buffer(440) := X"0C0007E2";
		ram_buffer(441) := X"00000000";
		ram_buffer(442) := X"AFA20010";
		ram_buffer(443) := X"27A40010";
		ram_buffer(444) := X"0C000CF0";
		ram_buffer(445) := X"24050002";
		ram_buffer(446) := X"8F848060";
		ram_buffer(447) := X"00003825";
		ram_buffer(448) := X"00003025";
		ram_buffer(449) := X"0C0003A3";
		ram_buffer(450) := X"00002825";
		ram_buffer(451) := X"1000FFF8";
		ram_buffer(452) := X"27A40010";
		ram_buffer(453) := X"27BDFFD0";
		ram_buffer(454) := X"AFB10020";
		ram_buffer(455) := X"3C110000";
		ram_buffer(456) := X"AFB30028";
		ram_buffer(457) := X"AFB20024";
		ram_buffer(458) := X"AFB0001C";
		ram_buffer(459) := X"AFBF002C";
		ram_buffer(460) := X"00008025";
		ram_buffer(461) := X"00009825";
		ram_buffer(462) := X"24120001";
		ram_buffer(463) := X"26316994";
		ram_buffer(464) := X"8F848064";
		ram_buffer(465) := X"00003825";
		ram_buffer(466) := X"00003025";
		ram_buffer(467) := X"0C000519";
		ram_buffer(468) := X"27A50010";
		ram_buffer(469) := X"1452000E";
		ram_buffer(470) := X"00001025";
		ram_buffer(471) := X"8FB30010";
		ram_buffer(472) := X"00000000";
		ram_buffer(473) := X"00132827";
		ram_buffer(474) := X"24040010";
		ram_buffer(475) := X"00521804";
		ram_buffer(476) := X"00651824";
		ram_buffer(477) := X"10600003";
		ram_buffer(478) := X"00021880";
		ram_buffer(479) := X"00711821";
		ram_buffer(480) := X"AC600000";
		ram_buffer(481) := X"24420001";
		ram_buffer(482) := X"1444FFF9";
		ram_buffer(483) := X"00521804";
		ram_buffer(484) := X"8F848060";
		ram_buffer(485) := X"00003825";
		ram_buffer(486) := X"00003025";
		ram_buffer(487) := X"0C000519";
		ram_buffer(488) := X"00002825";
		ram_buffer(489) := X"1452FFE6";
		ram_buffer(490) := X"00002025";
		ram_buffer(491) := X"240600F9";
		ram_buffer(492) := X"24050010";
		ram_buffer(493) := X"00921004";
		ram_buffer(494) := X"02621824";
		ram_buffer(495) := X"1060000A";
		ram_buffer(496) := X"00041880";
		ram_buffer(497) := X"00711821";
		ram_buffer(498) := X"8C670000";
		ram_buffer(499) := X"00000000";
		ram_buffer(500) := X"14E60011";
		ram_buffer(501) := X"00000000";
		ram_buffer(502) := X"AC600000";
		ram_buffer(503) := X"00501824";
		ram_buffer(504) := X"10600004";
		ram_buffer(505) := X"00000000";
		ram_buffer(506) := X"00021027";
		ram_buffer(507) := X"10000002";
		ram_buffer(508) := X"02028024";
		ram_buffer(509) := X"02028025";
		ram_buffer(510) := X"24840001";
		ram_buffer(511) := X"1485FFEE";
		ram_buffer(512) := X"00921004";
		ram_buffer(513) := X"8F82805C";
		ram_buffer(514) := X"00000000";
		ram_buffer(515) := X"AC500008";
		ram_buffer(516) := X"1000FFCB";
		ram_buffer(517) := X"00000000";
		ram_buffer(518) := X"8C620000";
		ram_buffer(519) := X"00000000";
		ram_buffer(520) := X"24420001";
		ram_buffer(521) := X"AC620000";
		ram_buffer(522) := X"1000FFF4";
		ram_buffer(523) := X"24840001";
		ram_buffer(524) := X"3C030000";
		ram_buffer(525) := X"8C626950";
		ram_buffer(526) := X"27BDFFE0";
		ram_buffer(527) := X"8C420004";
		ram_buffer(528) := X"AFB10018";
		ram_buffer(529) := X"3C110000";
		ram_buffer(530) := X"AFB00014";
		ram_buffer(531) := X"AFBF001C";
		ram_buffer(532) := X"00608025";
		ram_buffer(533) := X"26316954";
		ram_buffer(534) := X"2C430008";
		ram_buffer(535) := X"1460000C";
		ram_buffer(536) := X"000210C0";
		ram_buffer(537) := X"8F828048";
		ram_buffer(538) := X"00000000";
		ram_buffer(539) := X"10400012";
		ram_buffer(540) := X"00000000";
		ram_buffer(541) := X"8FBF001C";
		ram_buffer(542) := X"8FB10018";
		ram_buffer(543) := X"8FB00014";
		ram_buffer(544) := X"27BD0020";
		ram_buffer(545) := X"AF808048";
		ram_buffer(546) := X"08000883";
		ram_buffer(547) := X"00000000";
		ram_buffer(548) := X"02221021";
		ram_buffer(549) := X"8C430000";
		ram_buffer(550) := X"8C440004";
		ram_buffer(551) := X"0060F809";
		ram_buffer(552) := X"00000000";
		ram_buffer(553) := X"8E026950";
		ram_buffer(554) := X"00000000";
		ram_buffer(555) := X"8C420004";
		ram_buffer(556) := X"1000FFEA";
		ram_buffer(557) := X"2C430008";
		ram_buffer(558) := X"8FBF001C";
		ram_buffer(559) := X"8FB10018";
		ram_buffer(560) := X"8FB00014";
		ram_buffer(561) := X"03E00008";
		ram_buffer(562) := X"27BD0020";
		ram_buffer(563) := X"3C020000";
		ram_buffer(564) := X"8C426950";
		ram_buffer(565) := X"240300FF";
		ram_buffer(566) := X"03E00008";
		ram_buffer(567) := X"AC430000";
		ram_buffer(568) := X"3C020000";
		ram_buffer(569) := X"8C426950";
		ram_buffer(570) := X"00000000";
		ram_buffer(571) := X"03E00008";
		ram_buffer(572) := X"AC400000";
		ram_buffer(573) := X"8F82805C";
		ram_buffer(574) := X"00000000";
		ram_buffer(575) := X"AC450008";
		ram_buffer(576) := X"1000FFFF";
		ram_buffer(577) := X"00000000";
		ram_buffer(578) := X"10C0000D";
		ram_buffer(579) := X"00C53021";
		ram_buffer(580) := X"2402FFE0";
		ram_buffer(581) := X"00C21824";
		ram_buffer(582) := X"0066302B";
		ram_buffer(583) := X"00A22824";
		ram_buffer(584) := X"00063140";
		ram_buffer(585) := X"24620020";
		ram_buffer(586) := X"00463021";
		ram_buffer(587) := X"3C021000";
		ram_buffer(588) := X"00822021";
		ram_buffer(589) := X"2402FFE0";
		ram_buffer(590) := X"14C50003";
		ram_buffer(591) := X"00A21824";
		ram_buffer(592) := X"03E00008";
		ram_buffer(593) := X"00000000";
		ram_buffer(594) := X"AC830000";
		ram_buffer(595) := X"AC600000";
		ram_buffer(596) := X"1000FFF9";
		ram_buffer(597) := X"24A50020";
		ram_buffer(598) := X"24820008";
		ram_buffer(599) := X"2403FFFF";
		ram_buffer(600) := X"AC820004";
		ram_buffer(601) := X"AC830008";
		ram_buffer(602) := X"AC82000C";
		ram_buffer(603) := X"AC820010";
		ram_buffer(604) := X"03E00008";
		ram_buffer(605) := X"AC800000";
		ram_buffer(606) := X"03E00008";
		ram_buffer(607) := X"AC800010";
		ram_buffer(608) := X"8C820004";
		ram_buffer(609) := X"00000000";
		ram_buffer(610) := X"8C430008";
		ram_buffer(611) := X"ACA20004";
		ram_buffer(612) := X"ACA30008";
		ram_buffer(613) := X"8C430008";
		ram_buffer(614) := X"00000000";
		ram_buffer(615) := X"AC650004";
		ram_buffer(616) := X"AC450008";
		ram_buffer(617) := X"8C820000";
		ram_buffer(618) := X"ACA40010";
		ram_buffer(619) := X"24420001";
		ram_buffer(620) := X"03E00008";
		ram_buffer(621) := X"AC820000";
		ram_buffer(622) := X"8CA60000";
		ram_buffer(623) := X"2403FFFF";
		ram_buffer(624) := X"14C3000F";
		ram_buffer(625) := X"24820008";
		ram_buffer(626) := X"8C820010";
		ram_buffer(627) := X"00000000";
		ram_buffer(628) := X"8C430004";
		ram_buffer(629) := X"00000000";
		ram_buffer(630) := X"ACA30004";
		ram_buffer(631) := X"AC650008";
		ram_buffer(632) := X"ACA20008";
		ram_buffer(633) := X"AC450004";
		ram_buffer(634) := X"8C820000";
		ram_buffer(635) := X"ACA40010";
		ram_buffer(636) := X"24420001";
		ram_buffer(637) := X"03E00008";
		ram_buffer(638) := X"AC820000";
		ram_buffer(639) := X"00E01025";
		ram_buffer(640) := X"8C470004";
		ram_buffer(641) := X"00000000";
		ram_buffer(642) := X"8CE30000";
		ram_buffer(643) := X"00000000";
		ram_buffer(644) := X"00C3182B";
		ram_buffer(645) := X"1060FFF9";
		ram_buffer(646) := X"00000000";
		ram_buffer(647) := X"1000FFEC";
		ram_buffer(648) := X"00000000";
		ram_buffer(649) := X"8C850004";
		ram_buffer(650) := X"8C820008";
		ram_buffer(651) := X"8C830010";
		ram_buffer(652) := X"ACA20008";
		ram_buffer(653) := X"8C820008";
		ram_buffer(654) := X"00000000";
		ram_buffer(655) := X"AC450004";
		ram_buffer(656) := X"8C650004";
		ram_buffer(657) := X"00000000";
		ram_buffer(658) := X"14850002";
		ram_buffer(659) := X"00000000";
		ram_buffer(660) := X"AC620004";
		ram_buffer(661) := X"8C620000";
		ram_buffer(662) := X"AC800010";
		ram_buffer(663) := X"2442FFFF";
		ram_buffer(664) := X"03E00008";
		ram_buffer(665) := X"AC620000";
		ram_buffer(666) := X"27BDFFE0";
		ram_buffer(667) := X"AFB20018";
		ram_buffer(668) := X"00C09025";
		ram_buffer(669) := X"8C860040";
		ram_buffer(670) := X"AFB10014";
		ram_buffer(671) := X"AFB00010";
		ram_buffer(672) := X"AFBF001C";
		ram_buffer(673) := X"00808025";
		ram_buffer(674) := X"8C910038";
		ram_buffer(675) := X"14C00011";
		ram_buffer(676) := X"00000000";
		ram_buffer(677) := X"8C830000";
		ram_buffer(678) := X"00000000";
		ram_buffer(679) := X"14600005";
		ram_buffer(680) := X"00001025";
		ram_buffer(681) := X"8C840004";
		ram_buffer(682) := X"0C0009DC";
		ram_buffer(683) := X"00000000";
		ram_buffer(684) := X"AE000004";
		ram_buffer(685) := X"8FBF001C";
		ram_buffer(686) := X"26310001";
		ram_buffer(687) := X"AE110038";
		ram_buffer(688) := X"8FB20018";
		ram_buffer(689) := X"8FB10014";
		ram_buffer(690) := X"8FB00010";
		ram_buffer(691) := X"03E00008";
		ram_buffer(692) := X"27BD0020";
		ram_buffer(693) := X"16400010";
		ram_buffer(694) := X"00000000";
		ram_buffer(695) := X"8C840008";
		ram_buffer(696) := X"0C00103D";
		ram_buffer(697) := X"00000000";
		ram_buffer(698) := X"8E020008";
		ram_buffer(699) := X"8E030040";
		ram_buffer(700) := X"00000000";
		ram_buffer(701) := X"00431021";
		ram_buffer(702) := X"8E030004";
		ram_buffer(703) := X"AE020008";
		ram_buffer(704) := X"0043182B";
		ram_buffer(705) := X"1460FFEB";
		ram_buffer(706) := X"00001025";
		ram_buffer(707) := X"8E030000";
		ram_buffer(708) := X"1000FFE8";
		ram_buffer(709) := X"AE030008";
		ram_buffer(710) := X"8C84000C";
		ram_buffer(711) := X"0C00103D";
		ram_buffer(712) := X"00000000";
		ram_buffer(713) := X"8E030040";
		ram_buffer(714) := X"8E02000C";
		ram_buffer(715) := X"00031823";
		ram_buffer(716) := X"8E040000";
		ram_buffer(717) := X"00431021";
		ram_buffer(718) := X"AE02000C";
		ram_buffer(719) := X"0044102B";
		ram_buffer(720) := X"10400005";
		ram_buffer(721) := X"00000000";
		ram_buffer(722) := X"8E020004";
		ram_buffer(723) := X"00000000";
		ram_buffer(724) := X"00431821";
		ram_buffer(725) := X"AE03000C";
		ram_buffer(726) := X"24030002";
		ram_buffer(727) := X"1643FFD5";
		ram_buffer(728) := X"00001025";
		ram_buffer(729) := X"0011182B";
		ram_buffer(730) := X"1000FFD2";
		ram_buffer(731) := X"02238823";
		ram_buffer(732) := X"00801025";
		ram_buffer(733) := X"8C460040";
		ram_buffer(734) := X"00000000";
		ram_buffer(735) := X"10C0000E";
		ram_buffer(736) := X"00A02025";
		ram_buffer(737) := X"8C43000C";
		ram_buffer(738) := X"8C450004";
		ram_buffer(739) := X"00661821";
		ram_buffer(740) := X"AC43000C";
		ram_buffer(741) := X"0065182B";
		ram_buffer(742) := X"14600004";
		ram_buffer(743) := X"00000000";
		ram_buffer(744) := X"8C430000";
		ram_buffer(745) := X"00000000";
		ram_buffer(746) := X"AC43000C";
		ram_buffer(747) := X"8C45000C";
		ram_buffer(748) := X"0800103D";
		ram_buffer(749) := X"00000000";
		ram_buffer(750) := X"03E00008";
		ram_buffer(751) := X"00000000";
		ram_buffer(752) := X"27BDFFE0";
		ram_buffer(753) := X"AFB00010";
		ram_buffer(754) := X"AFB20018";
		ram_buffer(755) := X"AFB10014";
		ram_buffer(756) := X"AFBF001C";
		ram_buffer(757) := X"0C000A17";
		ram_buffer(758) := X"00808025";
		ram_buffer(759) := X"92110045";
		ram_buffer(760) := X"26120024";
		ram_buffer(761) := X"00118E00";
		ram_buffer(762) := X"00118E03";
		ram_buffer(763) := X"1E200013";
		ram_buffer(764) := X"2402FFFF";
		ram_buffer(765) := X"A2020045";
		ram_buffer(766) := X"0C000A2A";
		ram_buffer(767) := X"00000000";
		ram_buffer(768) := X"0C000A17";
		ram_buffer(769) := X"00000000";
		ram_buffer(770) := X"92110044";
		ram_buffer(771) := X"26120010";
		ram_buffer(772) := X"00118E00";
		ram_buffer(773) := X"00118E03";
		ram_buffer(774) := X"1E200016";
		ram_buffer(775) := X"2402FFFF";
		ram_buffer(776) := X"8FBF001C";
		ram_buffer(777) := X"8FB20018";
		ram_buffer(778) := X"8FB10014";
		ram_buffer(779) := X"A2020044";
		ram_buffer(780) := X"8FB00010";
		ram_buffer(781) := X"08000A2A";
		ram_buffer(782) := X"27BD0020";
		ram_buffer(783) := X"8E020024";
		ram_buffer(784) := X"00000000";
		ram_buffer(785) := X"1040FFEB";
		ram_buffer(786) := X"2402FFFF";
		ram_buffer(787) := X"0C0008FA";
		ram_buffer(788) := X"02402025";
		ram_buffer(789) := X"10400003";
		ram_buffer(790) := X"00000000";
		ram_buffer(791) := X"0C00097A";
		ram_buffer(792) := X"00000000";
		ram_buffer(793) := X"2631FFFF";
		ram_buffer(794) := X"00118E00";
		ram_buffer(795) := X"1000FFDF";
		ram_buffer(796) := X"00118E03";
		ram_buffer(797) := X"8E020010";
		ram_buffer(798) := X"00000000";
		ram_buffer(799) := X"1040FFE8";
		ram_buffer(800) := X"2402FFFF";
		ram_buffer(801) := X"0C0008FA";
		ram_buffer(802) := X"02402025";
		ram_buffer(803) := X"10400003";
		ram_buffer(804) := X"00000000";
		ram_buffer(805) := X"0C00097A";
		ram_buffer(806) := X"00000000";
		ram_buffer(807) := X"2631FFFF";
		ram_buffer(808) := X"00118E00";
		ram_buffer(809) := X"1000FFDC";
		ram_buffer(810) := X"00118E03";
		ram_buffer(811) := X"27BDFFE0";
		ram_buffer(812) := X"AFB10018";
		ram_buffer(813) := X"AFB00014";
		ram_buffer(814) := X"AFBF001C";
		ram_buffer(815) := X"00808025";
		ram_buffer(816) := X"14800005";
		ram_buffer(817) := X"00A08825";
		ram_buffer(818) := X"3C040000";
		ram_buffer(819) := X"2405011B";
		ram_buffer(820) := X"0C00023D";
		ram_buffer(821) := X"248445B4";
		ram_buffer(822) := X"0C000A17";
		ram_buffer(823) := X"00000000";
		ram_buffer(824) := X"8E050040";
		ram_buffer(825) := X"8E03003C";
		ram_buffer(826) := X"8E040000";
		ram_buffer(827) := X"00A30018";
		ram_buffer(828) := X"AE000038";
		ram_buffer(829) := X"AE040008";
		ram_buffer(830) := X"00001012";
		ram_buffer(831) := X"00821821";
		ram_buffer(832) := X"00451023";
		ram_buffer(833) := X"00821021";
		ram_buffer(834) := X"AE02000C";
		ram_buffer(835) := X"2402FFFF";
		ram_buffer(836) := X"A2020044";
		ram_buffer(837) := X"AE030004";
		ram_buffer(838) := X"A2020045";
		ram_buffer(839) := X"16200013";
		ram_buffer(840) := X"00000000";
		ram_buffer(841) := X"8E020010";
		ram_buffer(842) := X"00000000";
		ram_buffer(843) := X"10400007";
		ram_buffer(844) := X"00000000";
		ram_buffer(845) := X"0C0008FA";
		ram_buffer(846) := X"26040010";
		ram_buffer(847) := X"10400003";
		ram_buffer(848) := X"00000000";
		ram_buffer(849) := X"0C00017D";
		ram_buffer(850) := X"00000000";
		ram_buffer(851) := X"0C000A2A";
		ram_buffer(852) := X"00000000";
		ram_buffer(853) := X"8FBF001C";
		ram_buffer(854) := X"8FB10018";
		ram_buffer(855) := X"8FB00014";
		ram_buffer(856) := X"24020001";
		ram_buffer(857) := X"03E00008";
		ram_buffer(858) := X"27BD0020";
		ram_buffer(859) := X"0C000256";
		ram_buffer(860) := X"26040010";
		ram_buffer(861) := X"0C000256";
		ram_buffer(862) := X"26040024";
		ram_buffer(863) := X"1000FFF3";
		ram_buffer(864) := X"00000000";
		ram_buffer(865) := X"27BDFFE0";
		ram_buffer(866) := X"AFB20018";
		ram_buffer(867) := X"AFB10014";
		ram_buffer(868) := X"AFBF001C";
		ram_buffer(869) := X"AFB00010";
		ram_buffer(870) := X"00809025";
		ram_buffer(871) := X"14800005";
		ram_buffer(872) := X"00A08825";
		ram_buffer(873) := X"3C040000";
		ram_buffer(874) := X"24050188";
		ram_buffer(875) := X"0C00023D";
		ram_buffer(876) := X"248445B4";
		ram_buffer(877) := X"02510018";
		ram_buffer(878) := X"00002012";
		ram_buffer(879) := X"0C001008";
		ram_buffer(880) := X"24840048";
		ram_buffer(881) := X"10400009";
		ram_buffer(882) := X"00408025";
		ram_buffer(883) := X"1620000E";
		ram_buffer(884) := X"00000000";
		ram_buffer(885) := X"AE020000";
		ram_buffer(886) := X"AE12003C";
		ram_buffer(887) := X"AE110040";
		ram_buffer(888) := X"24050001";
		ram_buffer(889) := X"0C00032B";
		ram_buffer(890) := X"02002025";
		ram_buffer(891) := X"8FBF001C";
		ram_buffer(892) := X"02001025";
		ram_buffer(893) := X"8FB20018";
		ram_buffer(894) := X"8FB10014";
		ram_buffer(895) := X"8FB00010";
		ram_buffer(896) := X"03E00008";
		ram_buffer(897) := X"27BD0020";
		ram_buffer(898) := X"24420048";
		ram_buffer(899) := X"1000FFF2";
		ram_buffer(900) := X"AE020000";
		ram_buffer(901) := X"27BDFFE0";
		ram_buffer(902) := X"AFB10018";
		ram_buffer(903) := X"AFB00014";
		ram_buffer(904) := X"AFBF001C";
		ram_buffer(905) := X"00808025";
		ram_buffer(906) := X"14800005";
		ram_buffer(907) := X"00A08825";
		ram_buffer(908) := X"3C040000";
		ram_buffer(909) := X"240502BD";
		ram_buffer(910) := X"0C00023D";
		ram_buffer(911) := X"248445B4";
		ram_buffer(912) := X"0211102B";
		ram_buffer(913) := X"10400006";
		ram_buffer(914) := X"24060002";
		ram_buffer(915) := X"3C040000";
		ram_buffer(916) := X"240502BE";
		ram_buffer(917) := X"0C00023D";
		ram_buffer(918) := X"248445B4";
		ram_buffer(919) := X"24060002";
		ram_buffer(920) := X"00002825";
		ram_buffer(921) := X"0C000361";
		ram_buffer(922) := X"02002025";
		ram_buffer(923) := X"10400002";
		ram_buffer(924) := X"00000000";
		ram_buffer(925) := X"AC510038";
		ram_buffer(926) := X"8FBF001C";
		ram_buffer(927) := X"8FB10018";
		ram_buffer(928) := X"8FB00014";
		ram_buffer(929) := X"03E00008";
		ram_buffer(930) := X"27BD0020";
		ram_buffer(931) := X"27BDFFC0";
		ram_buffer(932) := X"AFB30028";
		ram_buffer(933) := X"AFB10020";
		ram_buffer(934) := X"AFB0001C";
		ram_buffer(935) := X"AFBF003C";
		ram_buffer(936) := X"AFB70038";
		ram_buffer(937) := X"AFB60034";
		ram_buffer(938) := X"AFB50030";
		ram_buffer(939) := X"AFB4002C";
		ram_buffer(940) := X"AFB20024";
		ram_buffer(941) := X"00808025";
		ram_buffer(942) := X"00A09825";
		ram_buffer(943) := X"AFA60048";
		ram_buffer(944) := X"14800005";
		ram_buffer(945) := X"00E08825";
		ram_buffer(946) := X"3C040000";
		ram_buffer(947) := X"240502D9";
		ram_buffer(948) := X"0C00023D";
		ram_buffer(949) := X"248445B4";
		ram_buffer(950) := X"16600006";
		ram_buffer(951) := X"24020002";
		ram_buffer(952) := X"8E020040";
		ram_buffer(953) := X"00000000";
		ram_buffer(954) := X"14400083";
		ram_buffer(955) := X"240502DA";
		ram_buffer(956) := X"24020002";
		ram_buffer(957) := X"16220005";
		ram_buffer(958) := X"24020001";
		ram_buffer(959) := X"8E03003C";
		ram_buffer(960) := X"00000000";
		ram_buffer(961) := X"14620081";
		ram_buffer(962) := X"3C040000";
		ram_buffer(963) := X"0C000991";
		ram_buffer(964) := X"00000000";
		ram_buffer(965) := X"14400009";
		ram_buffer(966) := X"0000B025";
		ram_buffer(967) := X"8FA20048";
		ram_buffer(968) := X"00000000";
		ram_buffer(969) := X"10400005";
		ram_buffer(970) := X"3C040000";
		ram_buffer(971) := X"240502DE";
		ram_buffer(972) := X"0C00023D";
		ram_buffer(973) := X"248445B4";
		ram_buffer(974) := X"0000B025";
		ram_buffer(975) := X"24150002";
		ram_buffer(976) := X"2412FFFF";
		ram_buffer(977) := X"1000003B";
		ram_buffer(978) := X"26140010";
		ram_buffer(979) := X"8FA20048";
		ram_buffer(980) := X"00000000";
		ram_buffer(981) := X"14400005";
		ram_buffer(982) := X"00000000";
		ram_buffer(983) := X"0C000A2A";
		ram_buffer(984) := X"00000000";
		ram_buffer(985) := X"1000004D";
		ram_buffer(986) := X"00001025";
		ram_buffer(987) := X"16C00003";
		ram_buffer(988) := X"00000000";
		ram_buffer(989) := X"0C000968";
		ram_buffer(990) := X"27A40010";
		ram_buffer(991) := X"0C000A2A";
		ram_buffer(992) := X"00000000";
		ram_buffer(993) := X"0C0007DC";
		ram_buffer(994) := X"00000000";
		ram_buffer(995) := X"0C000A17";
		ram_buffer(996) := X"00000000";
		ram_buffer(997) := X"92020044";
		ram_buffer(998) := X"00000000";
		ram_buffer(999) := X"00021600";
		ram_buffer(1000) := X"00021603";
		ram_buffer(1001) := X"14520002";
		ram_buffer(1002) := X"00000000";
		ram_buffer(1003) := X"A2000044";
		ram_buffer(1004) := X"92020045";
		ram_buffer(1005) := X"00000000";
		ram_buffer(1006) := X"00021600";
		ram_buffer(1007) := X"00021603";
		ram_buffer(1008) := X"14520002";
		ram_buffer(1009) := X"00000000";
		ram_buffer(1010) := X"A2000045";
		ram_buffer(1011) := X"0C000A2A";
		ram_buffer(1012) := X"00000000";
		ram_buffer(1013) := X"27A50048";
		ram_buffer(1014) := X"0C000DF0";
		ram_buffer(1015) := X"27A40010";
		ram_buffer(1016) := X"1440003F";
		ram_buffer(1017) := X"00000000";
		ram_buffer(1018) := X"0C000A17";
		ram_buffer(1019) := X"00000000";
		ram_buffer(1020) := X"8E170038";
		ram_buffer(1021) := X"8E16003C";
		ram_buffer(1022) := X"0C000A2A";
		ram_buffer(1023) := X"00000000";
		ram_buffer(1024) := X"16F60031";
		ram_buffer(1025) := X"00000000";
		ram_buffer(1026) := X"8FA50048";
		ram_buffer(1027) := X"0C0008C0";
		ram_buffer(1028) := X"02802025";
		ram_buffer(1029) := X"0C0002F0";
		ram_buffer(1030) := X"02002025";
		ram_buffer(1031) := X"0C000C85";
		ram_buffer(1032) := X"00000000";
		ram_buffer(1033) := X"14400003";
		ram_buffer(1034) := X"24160001";
		ram_buffer(1035) := X"0C00017D";
		ram_buffer(1036) := X"00000000";
		ram_buffer(1037) := X"0C000A17";
		ram_buffer(1038) := X"00000000";
		ram_buffer(1039) := X"8E020038";
		ram_buffer(1040) := X"8E03003C";
		ram_buffer(1041) := X"00000000";
		ram_buffer(1042) := X"0043102B";
		ram_buffer(1043) := X"14400003";
		ram_buffer(1044) := X"02203025";
		ram_buffer(1045) := X"1635FFBD";
		ram_buffer(1046) := X"00000000";
		ram_buffer(1047) := X"02602825";
		ram_buffer(1048) := X"0C00029A";
		ram_buffer(1049) := X"02002025";
		ram_buffer(1050) := X"8E030024";
		ram_buffer(1051) := X"00000000";
		ram_buffer(1052) := X"10600003";
		ram_buffer(1053) := X"00000000";
		ram_buffer(1054) := X"0C0008FA";
		ram_buffer(1055) := X"26040024";
		ram_buffer(1056) := X"10400003";
		ram_buffer(1057) := X"00000000";
		ram_buffer(1058) := X"0C00017D";
		ram_buffer(1059) := X"00000000";
		ram_buffer(1060) := X"0C000A2A";
		ram_buffer(1061) := X"00000000";
		ram_buffer(1062) := X"24020001";
		ram_buffer(1063) := X"8FBF003C";
		ram_buffer(1064) := X"8FB70038";
		ram_buffer(1065) := X"8FB60034";
		ram_buffer(1066) := X"8FB50030";
		ram_buffer(1067) := X"8FB4002C";
		ram_buffer(1068) := X"8FB30028";
		ram_buffer(1069) := X"8FB20024";
		ram_buffer(1070) := X"8FB10020";
		ram_buffer(1071) := X"8FB0001C";
		ram_buffer(1072) := X"03E00008";
		ram_buffer(1073) := X"27BD0040";
		ram_buffer(1074) := X"0C0002F0";
		ram_buffer(1075) := X"02002025";
		ram_buffer(1076) := X"0C000C85";
		ram_buffer(1077) := X"24160001";
		ram_buffer(1078) := X"1000FFD6";
		ram_buffer(1079) := X"00000000";
		ram_buffer(1080) := X"0C0002F0";
		ram_buffer(1081) := X"02002025";
		ram_buffer(1082) := X"0C000C85";
		ram_buffer(1083) := X"00000000";
		ram_buffer(1084) := X"1000FFEA";
		ram_buffer(1085) := X"00001025";
		ram_buffer(1086) := X"3C040000";
		ram_buffer(1087) := X"0C00023D";
		ram_buffer(1088) := X"248445B4";
		ram_buffer(1089) := X"1000FF7B";
		ram_buffer(1090) := X"24020002";
		ram_buffer(1091) := X"240502DB";
		ram_buffer(1092) := X"0C00023D";
		ram_buffer(1093) := X"248445B4";
		ram_buffer(1094) := X"1000FF7C";
		ram_buffer(1095) := X"00000000";
		ram_buffer(1096) := X"27BDFFE8";
		ram_buffer(1097) := X"00803025";
		ram_buffer(1098) := X"00002825";
		ram_buffer(1099) := X"AFB00010";
		ram_buffer(1100) := X"AFBF0014";
		ram_buffer(1101) := X"0C000361";
		ram_buffer(1102) := X"24040001";
		ram_buffer(1103) := X"10400009";
		ram_buffer(1104) := X"00408025";
		ram_buffer(1105) := X"AC400004";
		ram_buffer(1106) := X"AC400000";
		ram_buffer(1107) := X"AC40000C";
		ram_buffer(1108) := X"00003825";
		ram_buffer(1109) := X"00003025";
		ram_buffer(1110) := X"00002825";
		ram_buffer(1111) := X"0C0003A3";
		ram_buffer(1112) := X"00402025";
		ram_buffer(1113) := X"8FBF0014";
		ram_buffer(1114) := X"02001025";
		ram_buffer(1115) := X"8FB00010";
		ram_buffer(1116) := X"03E00008";
		ram_buffer(1117) := X"27BD0018";
		ram_buffer(1118) := X"27BDFFE0";
		ram_buffer(1119) := X"AFB00010";
		ram_buffer(1120) := X"AFBF001C";
		ram_buffer(1121) := X"AFB20018";
		ram_buffer(1122) := X"AFB10014";
		ram_buffer(1123) := X"14800005";
		ram_buffer(1124) := X"00808025";
		ram_buffer(1125) := X"3C040000";
		ram_buffer(1126) := X"24050241";
		ram_buffer(1127) := X"0C00023D";
		ram_buffer(1128) := X"248445B4";
		ram_buffer(1129) := X"8E120004";
		ram_buffer(1130) := X"0C00098E";
		ram_buffer(1131) := X"00008825";
		ram_buffer(1132) := X"1642000B";
		ram_buffer(1133) := X"00000000";
		ram_buffer(1134) := X"8E02000C";
		ram_buffer(1135) := X"24110001";
		ram_buffer(1136) := X"2442FFFF";
		ram_buffer(1137) := X"14400006";
		ram_buffer(1138) := X"AE02000C";
		ram_buffer(1139) := X"00003825";
		ram_buffer(1140) := X"00003025";
		ram_buffer(1141) := X"00002825";
		ram_buffer(1142) := X"0C0003A3";
		ram_buffer(1143) := X"02002025";
		ram_buffer(1144) := X"8FBF001C";
		ram_buffer(1145) := X"02201025";
		ram_buffer(1146) := X"8FB20018";
		ram_buffer(1147) := X"8FB10014";
		ram_buffer(1148) := X"8FB00010";
		ram_buffer(1149) := X"03E00008";
		ram_buffer(1150) := X"27BD0020";
		ram_buffer(1151) := X"27BDFFD0";
		ram_buffer(1152) := X"AFB40024";
		ram_buffer(1153) := X"AFB30020";
		ram_buffer(1154) := X"AFB2001C";
		ram_buffer(1155) := X"AFB00014";
		ram_buffer(1156) := X"AFBF002C";
		ram_buffer(1157) := X"AFB50028";
		ram_buffer(1158) := X"AFB10018";
		ram_buffer(1159) := X"00808025";
		ram_buffer(1160) := X"00A09825";
		ram_buffer(1161) := X"00C0A025";
		ram_buffer(1162) := X"14800005";
		ram_buffer(1163) := X"00E09025";
		ram_buffer(1164) := X"3C040000";
		ram_buffer(1165) := X"2405039F";
		ram_buffer(1166) := X"0C00023D";
		ram_buffer(1167) := X"248445B4";
		ram_buffer(1168) := X"16600006";
		ram_buffer(1169) := X"24020002";
		ram_buffer(1170) := X"8E020040";
		ram_buffer(1171) := X"00000000";
		ram_buffer(1172) := X"14400036";
		ram_buffer(1173) := X"240503A0";
		ram_buffer(1174) := X"24020002";
		ram_buffer(1175) := X"16420005";
		ram_buffer(1176) := X"24020001";
		ram_buffer(1177) := X"8E03003C";
		ram_buffer(1178) := X"00000000";
		ram_buffer(1179) := X"14620034";
		ram_buffer(1180) := X"240503A1";
		ram_buffer(1181) := X"8E020038";
		ram_buffer(1182) := X"8E03003C";
		ram_buffer(1183) := X"00000000";
		ram_buffer(1184) := X"0043102B";
		ram_buffer(1185) := X"14400003";
		ram_buffer(1186) := X"24030002";
		ram_buffer(1187) := X"16430018";
		ram_buffer(1188) := X"00000000";
		ram_buffer(1189) := X"92110045";
		ram_buffer(1190) := X"02403025";
		ram_buffer(1191) := X"0011AE00";
		ram_buffer(1192) := X"02602825";
		ram_buffer(1193) := X"0C00029A";
		ram_buffer(1194) := X"02002025";
		ram_buffer(1195) := X"0015AE03";
		ram_buffer(1196) := X"2402FFFF";
		ram_buffer(1197) := X"16A20017";
		ram_buffer(1198) := X"00000000";
		ram_buffer(1199) := X"8E020024";
		ram_buffer(1200) := X"00000000";
		ram_buffer(1201) := X"14400003";
		ram_buffer(1202) := X"00000000";
		ram_buffer(1203) := X"10000008";
		ram_buffer(1204) := X"24020001";
		ram_buffer(1205) := X"0C0008FA";
		ram_buffer(1206) := X"26040024";
		ram_buffer(1207) := X"1040FFFB";
		ram_buffer(1208) := X"00000000";
		ram_buffer(1209) := X"12800002";
		ram_buffer(1210) := X"24020001";
		ram_buffer(1211) := X"AE820000";
		ram_buffer(1212) := X"8FBF002C";
		ram_buffer(1213) := X"8FB50028";
		ram_buffer(1214) := X"8FB40024";
		ram_buffer(1215) := X"8FB30020";
		ram_buffer(1216) := X"8FB2001C";
		ram_buffer(1217) := X"8FB10018";
		ram_buffer(1218) := X"8FB00014";
		ram_buffer(1219) := X"03E00008";
		ram_buffer(1220) := X"27BD0030";
		ram_buffer(1221) := X"26310001";
		ram_buffer(1222) := X"00118E00";
		ram_buffer(1223) := X"00118E03";
		ram_buffer(1224) := X"A2110045";
		ram_buffer(1225) := X"1000FFF2";
		ram_buffer(1226) := X"24020001";
		ram_buffer(1227) := X"3C040000";
		ram_buffer(1228) := X"0C00023D";
		ram_buffer(1229) := X"248445B4";
		ram_buffer(1230) := X"1000FFC8";
		ram_buffer(1231) := X"24020002";
		ram_buffer(1232) := X"3C040000";
		ram_buffer(1233) := X"0C00023D";
		ram_buffer(1234) := X"248445B4";
		ram_buffer(1235) := X"1000FFC9";
		ram_buffer(1236) := X"00000000";
		ram_buffer(1237) := X"27BDFFE0";
		ram_buffer(1238) := X"AFB10018";
		ram_buffer(1239) := X"AFB00014";
		ram_buffer(1240) := X"AFBF001C";
		ram_buffer(1241) := X"00808025";
		ram_buffer(1242) := X"14800005";
		ram_buffer(1243) := X"00A08825";
		ram_buffer(1244) := X"3C040000";
		ram_buffer(1245) := X"2405043C";
		ram_buffer(1246) := X"0C00023D";
		ram_buffer(1247) := X"248445B4";
		ram_buffer(1248) := X"8E020040";
		ram_buffer(1249) := X"00000000";
		ram_buffer(1250) := X"10400004";
		ram_buffer(1251) := X"24050440";
		ram_buffer(1252) := X"3C040000";
		ram_buffer(1253) := X"0C00023D";
		ram_buffer(1254) := X"248445B4";
		ram_buffer(1255) := X"8E020000";
		ram_buffer(1256) := X"00000000";
		ram_buffer(1257) := X"14400005";
		ram_buffer(1258) := X"00000000";
		ram_buffer(1259) := X"8E020004";
		ram_buffer(1260) := X"00000000";
		ram_buffer(1261) := X"14400026";
		ram_buffer(1262) := X"3C040000";
		ram_buffer(1263) := X"8E030038";
		ram_buffer(1264) := X"8E04003C";
		ram_buffer(1265) := X"00000000";
		ram_buffer(1266) := X"0064202B";
		ram_buffer(1267) := X"10800016";
		ram_buffer(1268) := X"00001025";
		ram_buffer(1269) := X"92020045";
		ram_buffer(1270) := X"24630001";
		ram_buffer(1271) := X"00022600";
		ram_buffer(1272) := X"AE030038";
		ram_buffer(1273) := X"00042603";
		ram_buffer(1274) := X"2403FFFF";
		ram_buffer(1275) := X"14830013";
		ram_buffer(1276) := X"24420001";
		ram_buffer(1277) := X"8E020024";
		ram_buffer(1278) := X"00000000";
		ram_buffer(1279) := X"14400003";
		ram_buffer(1280) := X"00000000";
		ram_buffer(1281) := X"10000008";
		ram_buffer(1282) := X"24020001";
		ram_buffer(1283) := X"0C0008FA";
		ram_buffer(1284) := X"26040024";
		ram_buffer(1285) := X"1040FFFB";
		ram_buffer(1286) := X"00000000";
		ram_buffer(1287) := X"12200002";
		ram_buffer(1288) := X"24020001";
		ram_buffer(1289) := X"AE220000";
		ram_buffer(1290) := X"8FBF001C";
		ram_buffer(1291) := X"8FB10018";
		ram_buffer(1292) := X"8FB00014";
		ram_buffer(1293) := X"03E00008";
		ram_buffer(1294) := X"27BD0020";
		ram_buffer(1295) := X"00021600";
		ram_buffer(1296) := X"00021603";
		ram_buffer(1297) := X"A2020045";
		ram_buffer(1298) := X"1000FFF7";
		ram_buffer(1299) := X"24020001";
		ram_buffer(1300) := X"24050445";
		ram_buffer(1301) := X"0C00023D";
		ram_buffer(1302) := X"248445B4";
		ram_buffer(1303) := X"1000FFD7";
		ram_buffer(1304) := X"00000000";
		ram_buffer(1305) := X"27BDFFC8";
		ram_buffer(1306) := X"AFB5002C";
		ram_buffer(1307) := X"AFB30024";
		ram_buffer(1308) := X"AFB00018";
		ram_buffer(1309) := X"AFBF0034";
		ram_buffer(1310) := X"AFB60030";
		ram_buffer(1311) := X"AFB40028";
		ram_buffer(1312) := X"AFB20020";
		ram_buffer(1313) := X"AFB1001C";
		ram_buffer(1314) := X"00808025";
		ram_buffer(1315) := X"00A09825";
		ram_buffer(1316) := X"AFA60040";
		ram_buffer(1317) := X"14800005";
		ram_buffer(1318) := X"00E0A825";
		ram_buffer(1319) := X"3C040000";
		ram_buffer(1320) := X"240504DC";
		ram_buffer(1321) := X"0C00023D";
		ram_buffer(1322) := X"248445B4";
		ram_buffer(1323) := X"16600005";
		ram_buffer(1324) := X"00000000";
		ram_buffer(1325) := X"8E020040";
		ram_buffer(1326) := X"00000000";
		ram_buffer(1327) := X"14400096";
		ram_buffer(1328) := X"3C040000";
		ram_buffer(1329) := X"0C000991";
		ram_buffer(1330) := X"00000000";
		ram_buffer(1331) := X"14400009";
		ram_buffer(1332) := X"0000B025";
		ram_buffer(1333) := X"8FA20040";
		ram_buffer(1334) := X"00000000";
		ram_buffer(1335) := X"10400005";
		ram_buffer(1336) := X"3C040000";
		ram_buffer(1337) := X"240504E0";
		ram_buffer(1338) := X"0C00023D";
		ram_buffer(1339) := X"248445B4";
		ram_buffer(1340) := X"0000B025";
		ram_buffer(1341) := X"2412FFFF";
		ram_buffer(1342) := X"1000004B";
		ram_buffer(1343) := X"26140024";
		ram_buffer(1344) := X"8E020024";
		ram_buffer(1345) := X"AE12000C";
		ram_buffer(1346) := X"10400063";
		ram_buffer(1347) := X"26040024";
		ram_buffer(1348) := X"1000005B";
		ram_buffer(1349) := X"00000000";
		ram_buffer(1350) := X"8FA20040";
		ram_buffer(1351) := X"00000000";
		ram_buffer(1352) := X"14400005";
		ram_buffer(1353) := X"00000000";
		ram_buffer(1354) := X"0C000A2A";
		ram_buffer(1355) := X"00000000";
		ram_buffer(1356) := X"1000005C";
		ram_buffer(1357) := X"00001025";
		ram_buffer(1358) := X"16C00003";
		ram_buffer(1359) := X"00000000";
		ram_buffer(1360) := X"0C000968";
		ram_buffer(1361) := X"27A40010";
		ram_buffer(1362) := X"0C000A2A";
		ram_buffer(1363) := X"00000000";
		ram_buffer(1364) := X"0C0007DC";
		ram_buffer(1365) := X"00000000";
		ram_buffer(1366) := X"0C000A17";
		ram_buffer(1367) := X"00000000";
		ram_buffer(1368) := X"92020044";
		ram_buffer(1369) := X"00000000";
		ram_buffer(1370) := X"00021600";
		ram_buffer(1371) := X"00021603";
		ram_buffer(1372) := X"14520002";
		ram_buffer(1373) := X"00000000";
		ram_buffer(1374) := X"A2000044";
		ram_buffer(1375) := X"92020045";
		ram_buffer(1376) := X"00000000";
		ram_buffer(1377) := X"00021600";
		ram_buffer(1378) := X"00021603";
		ram_buffer(1379) := X"14520002";
		ram_buffer(1380) := X"00000000";
		ram_buffer(1381) := X"A2000045";
		ram_buffer(1382) := X"0C000A2A";
		ram_buffer(1383) := X"00000000";
		ram_buffer(1384) := X"27A50040";
		ram_buffer(1385) := X"0C000DF0";
		ram_buffer(1386) := X"27A40010";
		ram_buffer(1387) := X"1440004D";
		ram_buffer(1388) := X"00000000";
		ram_buffer(1389) := X"0C000A17";
		ram_buffer(1390) := X"00000000";
		ram_buffer(1391) := X"8E110038";
		ram_buffer(1392) := X"0C000A2A";
		ram_buffer(1393) := X"00000000";
		ram_buffer(1394) := X"16200040";
		ram_buffer(1395) := X"00000000";
		ram_buffer(1396) := X"8E020000";
		ram_buffer(1397) := X"00000000";
		ram_buffer(1398) := X"14400008";
		ram_buffer(1399) := X"00000000";
		ram_buffer(1400) := X"0C000A17";
		ram_buffer(1401) := X"00000000";
		ram_buffer(1402) := X"8E040004";
		ram_buffer(1403) := X"0C00099B";
		ram_buffer(1404) := X"00000000";
		ram_buffer(1405) := X"0C000A2A";
		ram_buffer(1406) := X"00000000";
		ram_buffer(1407) := X"8FA50040";
		ram_buffer(1408) := X"0C0008C0";
		ram_buffer(1409) := X"02802025";
		ram_buffer(1410) := X"0C0002F0";
		ram_buffer(1411) := X"02002025";
		ram_buffer(1412) := X"0C000C85";
		ram_buffer(1413) := X"00000000";
		ram_buffer(1414) := X"14400003";
		ram_buffer(1415) := X"24160001";
		ram_buffer(1416) := X"0C00017D";
		ram_buffer(1417) := X"00000000";
		ram_buffer(1418) := X"0C000A17";
		ram_buffer(1419) := X"00000000";
		ram_buffer(1420) := X"8E110038";
		ram_buffer(1421) := X"00000000";
		ram_buffer(1422) := X"1220FFB7";
		ram_buffer(1423) := X"02602825";
		ram_buffer(1424) := X"8E12000C";
		ram_buffer(1425) := X"0C0002DC";
		ram_buffer(1426) := X"02002025";
		ram_buffer(1427) := X"16A0FFAC";
		ram_buffer(1428) := X"2631FFFF";
		ram_buffer(1429) := X"8E020000";
		ram_buffer(1430) := X"AE110038";
		ram_buffer(1431) := X"14400004";
		ram_buffer(1432) := X"00000000";
		ram_buffer(1433) := X"0C000E35";
		ram_buffer(1434) := X"00000000";
		ram_buffer(1435) := X"AE020004";
		ram_buffer(1436) := X"8E020010";
		ram_buffer(1437) := X"00000000";
		ram_buffer(1438) := X"10400007";
		ram_buffer(1439) := X"26040010";
		ram_buffer(1440) := X"0C0008FA";
		ram_buffer(1441) := X"00000000";
		ram_buffer(1442) := X"10400003";
		ram_buffer(1443) := X"00000000";
		ram_buffer(1444) := X"0C00017D";
		ram_buffer(1445) := X"00000000";
		ram_buffer(1446) := X"0C000A2A";
		ram_buffer(1447) := X"00000000";
		ram_buffer(1448) := X"24020001";
		ram_buffer(1449) := X"8FBF0034";
		ram_buffer(1450) := X"8FB60030";
		ram_buffer(1451) := X"8FB5002C";
		ram_buffer(1452) := X"8FB40028";
		ram_buffer(1453) := X"8FB30024";
		ram_buffer(1454) := X"8FB20020";
		ram_buffer(1455) := X"8FB1001C";
		ram_buffer(1456) := X"8FB00018";
		ram_buffer(1457) := X"03E00008";
		ram_buffer(1458) := X"27BD0038";
		ram_buffer(1459) := X"0C0002F0";
		ram_buffer(1460) := X"02002025";
		ram_buffer(1461) := X"0C000C85";
		ram_buffer(1462) := X"24160001";
		ram_buffer(1463) := X"1000FFD2";
		ram_buffer(1464) := X"00000000";
		ram_buffer(1465) := X"0C0002F0";
		ram_buffer(1466) := X"02002025";
		ram_buffer(1467) := X"0C000C85";
		ram_buffer(1468) := X"00000000";
		ram_buffer(1469) := X"0C000A17";
		ram_buffer(1470) := X"00000000";
		ram_buffer(1471) := X"8E110038";
		ram_buffer(1472) := X"0C000A2A";
		ram_buffer(1473) := X"00000000";
		ram_buffer(1474) := X"1620FFC7";
		ram_buffer(1475) := X"24160001";
		ram_buffer(1476) := X"1000FFE4";
		ram_buffer(1477) := X"00001025";
		ram_buffer(1478) := X"240504DD";
		ram_buffer(1479) := X"0C00023D";
		ram_buffer(1480) := X"248445B4";
		ram_buffer(1481) := X"1000FF67";
		ram_buffer(1482) := X"00000000";
		ram_buffer(1483) := X"27BDFFE0";
		ram_buffer(1484) := X"AFB10014";
		ram_buffer(1485) := X"AFB00010";
		ram_buffer(1486) := X"AFBF001C";
		ram_buffer(1487) := X"AFB20018";
		ram_buffer(1488) := X"00808025";
		ram_buffer(1489) := X"14800005";
		ram_buffer(1490) := X"00A08825";
		ram_buffer(1491) := X"3C040000";
		ram_buffer(1492) := X"24050278";
		ram_buffer(1493) := X"0C00023D";
		ram_buffer(1494) := X"248445B4";
		ram_buffer(1495) := X"8E120004";
		ram_buffer(1496) := X"0C00098E";
		ram_buffer(1497) := X"00000000";
		ram_buffer(1498) := X"1642000C";
		ram_buffer(1499) := X"00003825";
		ram_buffer(1500) := X"8E02000C";
		ram_buffer(1501) := X"00000000";
		ram_buffer(1502) := X"24420001";
		ram_buffer(1503) := X"AE02000C";
		ram_buffer(1504) := X"24020001";
		ram_buffer(1505) := X"8FBF001C";
		ram_buffer(1506) := X"8FB20018";
		ram_buffer(1507) := X"8FB10014";
		ram_buffer(1508) := X"8FB00010";
		ram_buffer(1509) := X"03E00008";
		ram_buffer(1510) := X"27BD0020";
		ram_buffer(1511) := X"02203025";
		ram_buffer(1512) := X"00002825";
		ram_buffer(1513) := X"0C000519";
		ram_buffer(1514) := X"02002025";
		ram_buffer(1515) := X"1040FFF5";
		ram_buffer(1516) := X"00000000";
		ram_buffer(1517) := X"8E03000C";
		ram_buffer(1518) := X"00000000";
		ram_buffer(1519) := X"24630001";
		ram_buffer(1520) := X"1000FFF0";
		ram_buffer(1521) := X"AE03000C";
		ram_buffer(1522) := X"27BDFFD0";
		ram_buffer(1523) := X"AFB40024";
		ram_buffer(1524) := X"AFB30020";
		ram_buffer(1525) := X"AFB00014";
		ram_buffer(1526) := X"AFBF002C";
		ram_buffer(1527) := X"AFB50028";
		ram_buffer(1528) := X"AFB2001C";
		ram_buffer(1529) := X"AFB10018";
		ram_buffer(1530) := X"00808025";
		ram_buffer(1531) := X"00A09825";
		ram_buffer(1532) := X"14800005";
		ram_buffer(1533) := X"00C0A025";
		ram_buffer(1534) := X"3C040000";
		ram_buffer(1535) := X"240505A0";
		ram_buffer(1536) := X"0C00023D";
		ram_buffer(1537) := X"248445B4";
		ram_buffer(1538) := X"16600005";
		ram_buffer(1539) := X"00000000";
		ram_buffer(1540) := X"8E020040";
		ram_buffer(1541) := X"00000000";
		ram_buffer(1542) := X"1440002C";
		ram_buffer(1543) := X"240505A1";
		ram_buffer(1544) := X"8E120038";
		ram_buffer(1545) := X"00000000";
		ram_buffer(1546) := X"12400019";
		ram_buffer(1547) := X"00001025";
		ram_buffer(1548) := X"92110044";
		ram_buffer(1549) := X"02602825";
		ram_buffer(1550) := X"0011AE00";
		ram_buffer(1551) := X"0C0002DC";
		ram_buffer(1552) := X"02002025";
		ram_buffer(1553) := X"2652FFFF";
		ram_buffer(1554) := X"0015AE03";
		ram_buffer(1555) := X"2402FFFF";
		ram_buffer(1556) := X"AE120038";
		ram_buffer(1557) := X"16A20017";
		ram_buffer(1558) := X"00000000";
		ram_buffer(1559) := X"8E020010";
		ram_buffer(1560) := X"00000000";
		ram_buffer(1561) := X"14400003";
		ram_buffer(1562) := X"00000000";
		ram_buffer(1563) := X"10000008";
		ram_buffer(1564) := X"24020001";
		ram_buffer(1565) := X"0C0008FA";
		ram_buffer(1566) := X"26040010";
		ram_buffer(1567) := X"1040FFFB";
		ram_buffer(1568) := X"00000000";
		ram_buffer(1569) := X"12800002";
		ram_buffer(1570) := X"24020001";
		ram_buffer(1571) := X"AE820000";
		ram_buffer(1572) := X"8FBF002C";
		ram_buffer(1573) := X"8FB50028";
		ram_buffer(1574) := X"8FB40024";
		ram_buffer(1575) := X"8FB30020";
		ram_buffer(1576) := X"8FB2001C";
		ram_buffer(1577) := X"8FB10018";
		ram_buffer(1578) := X"8FB00014";
		ram_buffer(1579) := X"03E00008";
		ram_buffer(1580) := X"27BD0030";
		ram_buffer(1581) := X"26310001";
		ram_buffer(1582) := X"00118E00";
		ram_buffer(1583) := X"00118E03";
		ram_buffer(1584) := X"A2110044";
		ram_buffer(1585) := X"1000FFF2";
		ram_buffer(1586) := X"24020001";
		ram_buffer(1587) := X"3C040000";
		ram_buffer(1588) := X"0C00023D";
		ram_buffer(1589) := X"248445B4";
		ram_buffer(1590) := X"1000FFD1";
		ram_buffer(1591) := X"00000000";
		ram_buffer(1592) := X"27BDFFE0";
		ram_buffer(1593) := X"AFB10014";
		ram_buffer(1594) := X"AFB00010";
		ram_buffer(1595) := X"AFBF001C";
		ram_buffer(1596) := X"AFB20018";
		ram_buffer(1597) := X"00808025";
		ram_buffer(1598) := X"14800005";
		ram_buffer(1599) := X"00A08825";
		ram_buffer(1600) := X"3C040000";
		ram_buffer(1601) := X"240505FC";
		ram_buffer(1602) := X"0C00023D";
		ram_buffer(1603) := X"248445B4";
		ram_buffer(1604) := X"16200005";
		ram_buffer(1605) := X"00000000";
		ram_buffer(1606) := X"8E020040";
		ram_buffer(1607) := X"00000000";
		ram_buffer(1608) := X"14400018";
		ram_buffer(1609) := X"240505FD";
		ram_buffer(1610) := X"8E020040";
		ram_buffer(1611) := X"00000000";
		ram_buffer(1612) := X"14400004";
		ram_buffer(1613) := X"240505FE";
		ram_buffer(1614) := X"3C040000";
		ram_buffer(1615) := X"0C00023D";
		ram_buffer(1616) := X"248445B4";
		ram_buffer(1617) := X"8E030038";
		ram_buffer(1618) := X"00000000";
		ram_buffer(1619) := X"10600007";
		ram_buffer(1620) := X"00001025";
		ram_buffer(1621) := X"8E12000C";
		ram_buffer(1622) := X"02202825";
		ram_buffer(1623) := X"0C0002DC";
		ram_buffer(1624) := X"02002025";
		ram_buffer(1625) := X"AE12000C";
		ram_buffer(1626) := X"24020001";
		ram_buffer(1627) := X"8FBF001C";
		ram_buffer(1628) := X"8FB20018";
		ram_buffer(1629) := X"8FB10014";
		ram_buffer(1630) := X"8FB00010";
		ram_buffer(1631) := X"03E00008";
		ram_buffer(1632) := X"27BD0020";
		ram_buffer(1633) := X"3C040000";
		ram_buffer(1634) := X"0C00023D";
		ram_buffer(1635) := X"248445B4";
		ram_buffer(1636) := X"1000FFE5";
		ram_buffer(1637) := X"00000000";
		ram_buffer(1638) := X"27BDFFE8";
		ram_buffer(1639) := X"AFB00010";
		ram_buffer(1640) := X"AFBF0014";
		ram_buffer(1641) := X"14800005";
		ram_buffer(1642) := X"00808025";
		ram_buffer(1643) := X"3C040000";
		ram_buffer(1644) := X"2405062F";
		ram_buffer(1645) := X"0C00023D";
		ram_buffer(1646) := X"248445B4";
		ram_buffer(1647) := X"0C000A17";
		ram_buffer(1648) := X"00000000";
		ram_buffer(1649) := X"8E100038";
		ram_buffer(1650) := X"0C000A2A";
		ram_buffer(1651) := X"00000000";
		ram_buffer(1652) := X"8FBF0014";
		ram_buffer(1653) := X"02001025";
		ram_buffer(1654) := X"8FB00010";
		ram_buffer(1655) := X"03E00008";
		ram_buffer(1656) := X"27BD0018";
		ram_buffer(1657) := X"27BDFFE0";
		ram_buffer(1658) := X"AFB10018";
		ram_buffer(1659) := X"AFBF001C";
		ram_buffer(1660) := X"AFB00014";
		ram_buffer(1661) := X"14800005";
		ram_buffer(1662) := X"00808825";
		ram_buffer(1663) := X"3C040000";
		ram_buffer(1664) := X"24050641";
		ram_buffer(1665) := X"0C00023D";
		ram_buffer(1666) := X"248445B4";
		ram_buffer(1667) := X"0C000A17";
		ram_buffer(1668) := X"00000000";
		ram_buffer(1669) := X"8E220038";
		ram_buffer(1670) := X"8E30003C";
		ram_buffer(1671) := X"0C000A2A";
		ram_buffer(1672) := X"02028023";
		ram_buffer(1673) := X"8FBF001C";
		ram_buffer(1674) := X"02001025";
		ram_buffer(1675) := X"8FB10018";
		ram_buffer(1676) := X"8FB00014";
		ram_buffer(1677) := X"03E00008";
		ram_buffer(1678) := X"27BD0020";
		ram_buffer(1679) := X"27BDFFE8";
		ram_buffer(1680) := X"AFB00010";
		ram_buffer(1681) := X"AFBF0014";
		ram_buffer(1682) := X"14800005";
		ram_buffer(1683) := X"00808025";
		ram_buffer(1684) := X"3C040000";
		ram_buffer(1685) := X"24050651";
		ram_buffer(1686) := X"0C00023D";
		ram_buffer(1687) := X"248445B4";
		ram_buffer(1688) := X"8FBF0014";
		ram_buffer(1689) := X"8E020038";
		ram_buffer(1690) := X"8FB00010";
		ram_buffer(1691) := X"03E00008";
		ram_buffer(1692) := X"27BD0018";
		ram_buffer(1693) := X"27BDFFE8";
		ram_buffer(1694) := X"AFB00010";
		ram_buffer(1695) := X"AFBF0014";
		ram_buffer(1696) := X"14800005";
		ram_buffer(1697) := X"00808025";
		ram_buffer(1698) := X"3C040000";
		ram_buffer(1699) := X"24050793";
		ram_buffer(1700) := X"0C00023D";
		ram_buffer(1701) := X"248445B4";
		ram_buffer(1702) := X"8E020038";
		ram_buffer(1703) := X"8FBF0014";
		ram_buffer(1704) := X"8FB00010";
		ram_buffer(1705) := X"2C420001";
		ram_buffer(1706) := X"03E00008";
		ram_buffer(1707) := X"27BD0018";
		ram_buffer(1708) := X"27BDFFE8";
		ram_buffer(1709) := X"AFB00010";
		ram_buffer(1710) := X"AFBF0014";
		ram_buffer(1711) := X"14800005";
		ram_buffer(1712) := X"00808025";
		ram_buffer(1713) := X"3C040000";
		ram_buffer(1714) := X"240507BA";
		ram_buffer(1715) := X"0C00023D";
		ram_buffer(1716) := X"248445B4";
		ram_buffer(1717) := X"8E030038";
		ram_buffer(1718) := X"8E02003C";
		ram_buffer(1719) := X"8FBF0014";
		ram_buffer(1720) := X"00431026";
		ram_buffer(1721) := X"8FB00010";
		ram_buffer(1722) := X"2C420001";
		ram_buffer(1723) := X"03E00008";
		ram_buffer(1724) := X"27BD0018";
		ram_buffer(1725) := X"3C030000";
		ram_buffer(1726) := X"246369D4";
		ram_buffer(1727) := X"00001025";
		ram_buffer(1728) := X"00603025";
		ram_buffer(1729) := X"2407000A";
		ram_buffer(1730) := X"8C680000";
		ram_buffer(1731) := X"00000000";
		ram_buffer(1732) := X"15000007";
		ram_buffer(1733) := X"24420001";
		ram_buffer(1734) := X"2442FFFF";
		ram_buffer(1735) := X"000210C0";
		ram_buffer(1736) := X"00C21021";
		ram_buffer(1737) := X"AC450000";
		ram_buffer(1738) := X"03E00008";
		ram_buffer(1739) := X"AC440004";
		ram_buffer(1740) := X"1447FFF5";
		ram_buffer(1741) := X"24630008";
		ram_buffer(1742) := X"03E00008";
		ram_buffer(1743) := X"00000000";
		ram_buffer(1744) := X"3C030000";
		ram_buffer(1745) := X"246369D4";
		ram_buffer(1746) := X"00001025";
		ram_buffer(1747) := X"00602825";
		ram_buffer(1748) := X"2406000A";
		ram_buffer(1749) := X"8C670004";
		ram_buffer(1750) := X"00000000";
		ram_buffer(1751) := X"14E40007";
		ram_buffer(1752) := X"24420001";
		ram_buffer(1753) := X"2442FFFF";
		ram_buffer(1754) := X"000210C0";
		ram_buffer(1755) := X"00A21021";
		ram_buffer(1756) := X"8C420000";
		ram_buffer(1757) := X"03E00008";
		ram_buffer(1758) := X"00000000";
		ram_buffer(1759) := X"1446FFF5";
		ram_buffer(1760) := X"24630008";
		ram_buffer(1761) := X"03E00008";
		ram_buffer(1762) := X"00001025";
		ram_buffer(1763) := X"3C030000";
		ram_buffer(1764) := X"246369D4";
		ram_buffer(1765) := X"00001025";
		ram_buffer(1766) := X"00602825";
		ram_buffer(1767) := X"2406000A";
		ram_buffer(1768) := X"8C670004";
		ram_buffer(1769) := X"00000000";
		ram_buffer(1770) := X"14E40007";
		ram_buffer(1771) := X"24420001";
		ram_buffer(1772) := X"2442FFFF";
		ram_buffer(1773) := X"000210C0";
		ram_buffer(1774) := X"00A21021";
		ram_buffer(1775) := X"AC400000";
		ram_buffer(1776) := X"03E00008";
		ram_buffer(1777) := X"AC400004";
		ram_buffer(1778) := X"1446FFF5";
		ram_buffer(1779) := X"24630008";
		ram_buffer(1780) := X"03E00008";
		ram_buffer(1781) := X"00000000";
		ram_buffer(1782) := X"27BDFFE8";
		ram_buffer(1783) := X"AFB00010";
		ram_buffer(1784) := X"AFBF0014";
		ram_buffer(1785) := X"14800005";
		ram_buffer(1786) := X"00808025";
		ram_buffer(1787) := X"3C040000";
		ram_buffer(1788) := X"2405065D";
		ram_buffer(1789) := X"0C00023D";
		ram_buffer(1790) := X"248445B4";
		ram_buffer(1791) := X"0C0006E3";
		ram_buffer(1792) := X"02002025";
		ram_buffer(1793) := X"8FBF0014";
		ram_buffer(1794) := X"02002025";
		ram_buffer(1795) := X"8FB00010";
		ram_buffer(1796) := X"08001030";
		ram_buffer(1797) := X"27BD0018";
		ram_buffer(1798) := X"8C820000";
		ram_buffer(1799) := X"00000000";
		ram_buffer(1800) := X"10400027";
		ram_buffer(1801) := X"24870008";
		ram_buffer(1802) := X"8C820004";
		ram_buffer(1803) := X"00000000";
		ram_buffer(1804) := X"8C420004";
		ram_buffer(1805) := X"00000000";
		ram_buffer(1806) := X"14470004";
		ram_buffer(1807) := X"AC820004";
		ram_buffer(1808) := X"8C82000C";
		ram_buffer(1809) := X"00000000";
		ram_buffer(1810) := X"AC820004";
		ram_buffer(1811) := X"8C820004";
		ram_buffer(1812) := X"00000000";
		ram_buffer(1813) := X"8C49000C";
		ram_buffer(1814) := X"8C820004";
		ram_buffer(1815) := X"00000000";
		ram_buffer(1816) := X"8C420004";
		ram_buffer(1817) := X"00000000";
		ram_buffer(1818) := X"14E20004";
		ram_buffer(1819) := X"AC820004";
		ram_buffer(1820) := X"8C82000C";
		ram_buffer(1821) := X"00000000";
		ram_buffer(1822) := X"AC820004";
		ram_buffer(1823) := X"8C820004";
		ram_buffer(1824) := X"00A03025";
		ram_buffer(1825) := X"8C42000C";
		ram_buffer(1826) := X"00000000";
		ram_buffer(1827) := X"24430034";
		ram_buffer(1828) := X"244A0044";
		ram_buffer(1829) := X"806B0000";
		ram_buffer(1830) := X"80C80000";
		ram_buffer(1831) := X"00000000";
		ram_buffer(1832) := X"150B0005";
		ram_buffer(1833) := X"00000000";
		ram_buffer(1834) := X"11000006";
		ram_buffer(1835) := X"24630001";
		ram_buffer(1836) := X"146AFFF8";
		ram_buffer(1837) := X"24C60001";
		ram_buffer(1838) := X"1522FFE7";
		ram_buffer(1839) := X"00000000";
		ram_buffer(1840) := X"00001025";
		ram_buffer(1841) := X"03E00008";
		ram_buffer(1842) := X"00000000";
		ram_buffer(1843) := X"8F828044";
		ram_buffer(1844) := X"00000000";
		ram_buffer(1845) := X"8C420000";
		ram_buffer(1846) := X"00000000";
		ram_buffer(1847) := X"14400005";
		ram_buffer(1848) := X"00000000";
		ram_buffer(1849) := X"2402FFFF";
		ram_buffer(1850) := X"AF828018";
		ram_buffer(1851) := X"03E00008";
		ram_buffer(1852) := X"00000000";
		ram_buffer(1853) := X"8F828044";
		ram_buffer(1854) := X"00000000";
		ram_buffer(1855) := X"8C42000C";
		ram_buffer(1856) := X"00000000";
		ram_buffer(1857) := X"8C42000C";
		ram_buffer(1858) := X"00000000";
		ram_buffer(1859) := X"8C420004";
		ram_buffer(1860) := X"1000FFF5";
		ram_buffer(1861) := X"00000000";
		ram_buffer(1862) := X"27BDFFE8";
		ram_buffer(1863) := X"AFB00010";
		ram_buffer(1864) := X"AFBF0014";
		ram_buffer(1865) := X"14800005";
		ram_buffer(1866) := X"00808025";
		ram_buffer(1867) := X"3C040000";
		ram_buffer(1868) := X"24050688";
		ram_buffer(1869) := X"0C00023D";
		ram_buffer(1870) := X"248445CC";
		ram_buffer(1871) := X"3C030000";
		ram_buffer(1872) := X"8E040014";
		ram_buffer(1873) := X"24634680";
		ram_buffer(1874) := X"14830007";
		ram_buffer(1875) := X"00001025";
		ram_buffer(1876) := X"3C030000";
		ram_buffer(1877) := X"8E040028";
		ram_buffer(1878) := X"246346A8";
		ram_buffer(1879) := X"10830002";
		ram_buffer(1880) := X"00000000";
		ram_buffer(1881) := X"2C820001";
		ram_buffer(1882) := X"8FBF0014";
		ram_buffer(1883) := X"8FB00010";
		ram_buffer(1884) := X"03E00008";
		ram_buffer(1885) := X"27BD0018";
		ram_buffer(1886) := X"27BDFFE0";
		ram_buffer(1887) := X"AFB10014";
		ram_buffer(1888) := X"AFB00010";
		ram_buffer(1889) := X"8F918034";
		ram_buffer(1890) := X"00808025";
		ram_buffer(1891) := X"8F82800C";
		ram_buffer(1892) := X"8F84800C";
		ram_buffer(1893) := X"AFB20018";
		ram_buffer(1894) := X"AFBF001C";
		ram_buffer(1895) := X"24840004";
		ram_buffer(1896) := X"A0400055";
		ram_buffer(1897) := X"0C000289";
		ram_buffer(1898) := X"00A09025";
		ram_buffer(1899) := X"2402FFFF";
		ram_buffer(1900) := X"1602000D";
		ram_buffer(1901) := X"00000000";
		ram_buffer(1902) := X"1240000C";
		ram_buffer(1903) := X"02308021";
		ram_buffer(1904) := X"8F85800C";
		ram_buffer(1905) := X"8FBF001C";
		ram_buffer(1906) := X"8FB20018";
		ram_buffer(1907) := X"8FB10014";
		ram_buffer(1908) := X"8FB00010";
		ram_buffer(1909) := X"3C040000";
		ram_buffer(1910) := X"24A50004";
		ram_buffer(1911) := X"24844680";
		ram_buffer(1912) := X"08000260";
		ram_buffer(1913) := X"27BD0020";
		ram_buffer(1914) := X"02308021";
		ram_buffer(1915) := X"8F82800C";
		ram_buffer(1916) := X"0211882B";
		ram_buffer(1917) := X"1220000A";
		ram_buffer(1918) := X"AC500004";
		ram_buffer(1919) := X"8F848040";
		ram_buffer(1920) := X"8F85800C";
		ram_buffer(1921) := X"8FBF001C";
		ram_buffer(1922) := X"8FB20018";
		ram_buffer(1923) := X"8FB10014";
		ram_buffer(1924) := X"8FB00010";
		ram_buffer(1925) := X"24A50004";
		ram_buffer(1926) := X"0800026E";
		ram_buffer(1927) := X"27BD0020";
		ram_buffer(1928) := X"8F848044";
		ram_buffer(1929) := X"8F85800C";
		ram_buffer(1930) := X"0C00026E";
		ram_buffer(1931) := X"24A50004";
		ram_buffer(1932) := X"8F828018";
		ram_buffer(1933) := X"00000000";
		ram_buffer(1934) := X"0202102B";
		ram_buffer(1935) := X"10400002";
		ram_buffer(1936) := X"00000000";
		ram_buffer(1937) := X"AF908018";
		ram_buffer(1938) := X"8FBF001C";
		ram_buffer(1939) := X"8FB20018";
		ram_buffer(1940) := X"8FB10014";
		ram_buffer(1941) := X"8FB00010";
		ram_buffer(1942) := X"03E00008";
		ram_buffer(1943) := X"27BD0020";
		ram_buffer(1944) := X"14800003";
		ram_buffer(1945) := X"00000000";
		ram_buffer(1946) := X"8F84800C";
		ram_buffer(1947) := X"00000000";
		ram_buffer(1948) := X"8C82002C";
		ram_buffer(1949) := X"03E00008";
		ram_buffer(1950) := X"00000000";
		ram_buffer(1951) := X"27BDFFE0";
		ram_buffer(1952) := X"AFB10014";
		ram_buffer(1953) := X"AFBF001C";
		ram_buffer(1954) := X"AFB20018";
		ram_buffer(1955) := X"AFB00010";
		ram_buffer(1956) := X"14800005";
		ram_buffer(1957) := X"00808825";
		ram_buffer(1958) := X"3C040000";
		ram_buffer(1959) := X"240506E9";
		ram_buffer(1960) := X"0C00023D";
		ram_buffer(1961) := X"248445CC";
		ram_buffer(1962) := X"0C000746";
		ram_buffer(1963) := X"02202025";
		ram_buffer(1964) := X"1040001C";
		ram_buffer(1965) := X"00008025";
		ram_buffer(1966) := X"8F828010";
		ram_buffer(1967) := X"00000000";
		ram_buffer(1968) := X"1440001F";
		ram_buffer(1969) := X"3C040000";
		ram_buffer(1970) := X"8F82800C";
		ram_buffer(1971) := X"8E30002C";
		ram_buffer(1972) := X"8C42002C";
		ram_buffer(1973) := X"26320004";
		ram_buffer(1974) := X"02402025";
		ram_buffer(1975) := X"0C000289";
		ram_buffer(1976) := X"0202802B";
		ram_buffer(1977) := X"8E24002C";
		ram_buffer(1978) := X"8F828030";
		ram_buffer(1979) := X"00000000";
		ram_buffer(1980) := X"0044102B";
		ram_buffer(1981) := X"10400002";
		ram_buffer(1982) := X"3A100001";
		ram_buffer(1983) := X"AF848030";
		ram_buffer(1984) := X"00041080";
		ram_buffer(1985) := X"00441021";
		ram_buffer(1986) := X"3C040000";
		ram_buffer(1987) := X"00021080";
		ram_buffer(1988) := X"248446E4";
		ram_buffer(1989) := X"02402825";
		ram_buffer(1990) := X"00822021";
		ram_buffer(1991) := X"0C000260";
		ram_buffer(1992) := X"00000000";
		ram_buffer(1993) := X"8FBF001C";
		ram_buffer(1994) := X"02001025";
		ram_buffer(1995) := X"8FB20018";
		ram_buffer(1996) := X"8FB10014";
		ram_buffer(1997) := X"8FB00010";
		ram_buffer(1998) := X"03E00008";
		ram_buffer(1999) := X"27BD0020";
		ram_buffer(2000) := X"26250018";
		ram_buffer(2001) := X"1000FFF5";
		ram_buffer(2002) := X"248446A8";
		ram_buffer(2003) := X"27BDFFE8";
		ram_buffer(2004) := X"AFBF0014";
		ram_buffer(2005) := X"0C000238";
		ram_buffer(2006) := X"00000000";
		ram_buffer(2007) := X"8FBF0014";
		ram_buffer(2008) := X"27BD0018";
		ram_buffer(2009) := X"AF80802C";
		ram_buffer(2010) := X"08001004";
		ram_buffer(2011) := X"00000000";
		ram_buffer(2012) := X"8F828010";
		ram_buffer(2013) := X"00000000";
		ram_buffer(2014) := X"24420001";
		ram_buffer(2015) := X"AF828010";
		ram_buffer(2016) := X"03E00008";
		ram_buffer(2017) := X"00000000";
		ram_buffer(2018) := X"8F828034";
		ram_buffer(2019) := X"03E00008";
		ram_buffer(2020) := X"00000000";
		ram_buffer(2021) := X"8F828034";
		ram_buffer(2022) := X"03E00008";
		ram_buffer(2023) := X"00000000";
		ram_buffer(2024) := X"8F828038";
		ram_buffer(2025) := X"03E00008";
		ram_buffer(2026) := X"00000000";
		ram_buffer(2027) := X"27BDFFE8";
		ram_buffer(2028) := X"AFB00010";
		ram_buffer(2029) := X"AFBF0014";
		ram_buffer(2030) := X"14800008";
		ram_buffer(2031) := X"00808025";
		ram_buffer(2032) := X"8F90800C";
		ram_buffer(2033) := X"00000000";
		ram_buffer(2034) := X"16000004";
		ram_buffer(2035) := X"24050893";
		ram_buffer(2036) := X"3C040000";
		ram_buffer(2037) := X"0C00023D";
		ram_buffer(2038) := X"248445CC";
		ram_buffer(2039) := X"8FBF0014";
		ram_buffer(2040) := X"26020034";
		ram_buffer(2041) := X"8FB00010";
		ram_buffer(2042) := X"03E00008";
		ram_buffer(2043) := X"27BD0018";
		ram_buffer(2044) := X"8F828014";
		ram_buffer(2045) := X"27BDFFE8";
		ram_buffer(2046) := X"14400005";
		ram_buffer(2047) := X"AFBF0014";
		ram_buffer(2048) := X"3C040000";
		ram_buffer(2049) := X"24050966";
		ram_buffer(2050) := X"0C00023D";
		ram_buffer(2051) := X"248445CC";
		ram_buffer(2052) := X"8FBF0014";
		ram_buffer(2053) := X"8F828014";
		ram_buffer(2054) := X"03E00008";
		ram_buffer(2055) := X"27BD0018";
		ram_buffer(2056) := X"8F828010";
		ram_buffer(2057) := X"27BDFFD8";
		ram_buffer(2058) := X"AFBF0024";
		ram_buffer(2059) := X"AFB40020";
		ram_buffer(2060) := X"AFB3001C";
		ram_buffer(2061) := X"AFB20018";
		ram_buffer(2062) := X"AFB10014";
		ram_buffer(2063) := X"1440006D";
		ram_buffer(2064) := X"AFB00010";
		ram_buffer(2065) := X"8F918034";
		ram_buffer(2066) := X"00000000";
		ram_buffer(2067) := X"26310001";
		ram_buffer(2068) := X"AF918034";
		ram_buffer(2069) := X"16200015";
		ram_buffer(2070) := X"00000000";
		ram_buffer(2071) := X"8F828044";
		ram_buffer(2072) := X"00000000";
		ram_buffer(2073) := X"8C420000";
		ram_buffer(2074) := X"00000000";
		ram_buffer(2075) := X"10400004";
		ram_buffer(2076) := X"240509E4";
		ram_buffer(2077) := X"3C040000";
		ram_buffer(2078) := X"0C00023D";
		ram_buffer(2079) := X"248445CC";
		ram_buffer(2080) := X"8F828044";
		ram_buffer(2081) := X"8F838040";
		ram_buffer(2082) := X"00000000";
		ram_buffer(2083) := X"AF838044";
		ram_buffer(2084) := X"AF828040";
		ram_buffer(2085) := X"8F828020";
		ram_buffer(2086) := X"00000000";
		ram_buffer(2087) := X"24420001";
		ram_buffer(2088) := X"AF828020";
		ram_buffer(2089) := X"0C000733";
		ram_buffer(2090) := X"00000000";
		ram_buffer(2091) := X"8F828018";
		ram_buffer(2092) := X"3C100000";
		ram_buffer(2093) := X"0222102B";
		ram_buffer(2094) := X"261046E4";
		ram_buffer(2095) := X"14400008";
		ram_buffer(2096) := X"00009825";
		ram_buffer(2097) := X"8F828044";
		ram_buffer(2098) := X"00000000";
		ram_buffer(2099) := X"8C420000";
		ram_buffer(2100) := X"00000000";
		ram_buffer(2101) := X"1440001E";
		ram_buffer(2102) := X"2402FFFF";
		ram_buffer(2103) := X"AF828018";
		ram_buffer(2104) := X"8F82800C";
		ram_buffer(2105) := X"00000000";
		ram_buffer(2106) := X"8C43002C";
		ram_buffer(2107) := X"00000000";
		ram_buffer(2108) := X"00031080";
		ram_buffer(2109) := X"00431021";
		ram_buffer(2110) := X"00021080";
		ram_buffer(2111) := X"02028021";
		ram_buffer(2112) := X"8E020000";
		ram_buffer(2113) := X"00000000";
		ram_buffer(2114) := X"2C420002";
		ram_buffer(2115) := X"14400002";
		ram_buffer(2116) := X"00000000";
		ram_buffer(2117) := X"24130001";
		ram_buffer(2118) := X"8F828024";
		ram_buffer(2119) := X"00000000";
		ram_buffer(2120) := X"10400002";
		ram_buffer(2121) := X"00000000";
		ram_buffer(2122) := X"24130001";
		ram_buffer(2123) := X"8FBF0024";
		ram_buffer(2124) := X"02601025";
		ram_buffer(2125) := X"8FB40020";
		ram_buffer(2126) := X"8FB3001C";
		ram_buffer(2127) := X"8FB20018";
		ram_buffer(2128) := X"8FB10014";
		ram_buffer(2129) := X"8FB00010";
		ram_buffer(2130) := X"03E00008";
		ram_buffer(2131) := X"27BD0028";
		ram_buffer(2132) := X"8F828044";
		ram_buffer(2133) := X"00000000";
		ram_buffer(2134) := X"8C42000C";
		ram_buffer(2135) := X"00000000";
		ram_buffer(2136) := X"8C52000C";
		ram_buffer(2137) := X"00000000";
		ram_buffer(2138) := X"8E420004";
		ram_buffer(2139) := X"00000000";
		ram_buffer(2140) := X"0222182B";
		ram_buffer(2141) := X"1460FFD9";
		ram_buffer(2142) := X"26540004";
		ram_buffer(2143) := X"0C000289";
		ram_buffer(2144) := X"02802025";
		ram_buffer(2145) := X"8E420028";
		ram_buffer(2146) := X"00000000";
		ram_buffer(2147) := X"10400003";
		ram_buffer(2148) := X"00000000";
		ram_buffer(2149) := X"0C000289";
		ram_buffer(2150) := X"26440018";
		ram_buffer(2151) := X"8E42002C";
		ram_buffer(2152) := X"8F838030";
		ram_buffer(2153) := X"00000000";
		ram_buffer(2154) := X"0062182B";
		ram_buffer(2155) := X"10600002";
		ram_buffer(2156) := X"00000000";
		ram_buffer(2157) := X"AF828030";
		ram_buffer(2158) := X"00022080";
		ram_buffer(2159) := X"00822021";
		ram_buffer(2160) := X"00042080";
		ram_buffer(2161) := X"02802825";
		ram_buffer(2162) := X"0C000260";
		ram_buffer(2163) := X"02042021";
		ram_buffer(2164) := X"8F83800C";
		ram_buffer(2165) := X"8E42002C";
		ram_buffer(2166) := X"8C63002C";
		ram_buffer(2167) := X"00000000";
		ram_buffer(2168) := X"0043102B";
		ram_buffer(2169) := X"1440FFB7";
		ram_buffer(2170) := X"00000000";
		ram_buffer(2171) := X"1000FFB5";
		ram_buffer(2172) := X"24130001";
		ram_buffer(2173) := X"8F828028";
		ram_buffer(2174) := X"00009825";
		ram_buffer(2175) := X"24420001";
		ram_buffer(2176) := X"AF828028";
		ram_buffer(2177) := X"1000FFC4";
		ram_buffer(2178) := X"00000000";
		ram_buffer(2179) := X"8F828010";
		ram_buffer(2180) := X"27BDFFD8";
		ram_buffer(2181) := X"AFBF0024";
		ram_buffer(2182) := X"AFB30020";
		ram_buffer(2183) := X"AFB2001C";
		ram_buffer(2184) := X"AFB10018";
		ram_buffer(2185) := X"1040000A";
		ram_buffer(2186) := X"AFB00014";
		ram_buffer(2187) := X"24020001";
		ram_buffer(2188) := X"AF828024";
		ram_buffer(2189) := X"8FBF0024";
		ram_buffer(2190) := X"8FB30020";
		ram_buffer(2191) := X"8FB2001C";
		ram_buffer(2192) := X"8FB10018";
		ram_buffer(2193) := X"8FB00014";
		ram_buffer(2194) := X"03E00008";
		ram_buffer(2195) := X"27BD0028";
		ram_buffer(2196) := X"AF808024";
		ram_buffer(2197) := X"8F908030";
		ram_buffer(2198) := X"3C120000";
		ram_buffer(2199) := X"00108880";
		ram_buffer(2200) := X"02308821";
		ram_buffer(2201) := X"00118880";
		ram_buffer(2202) := X"265246E4";
		ram_buffer(2203) := X"3C130000";
		ram_buffer(2204) := X"02518821";
		ram_buffer(2205) := X"267345CC";
		ram_buffer(2206) := X"8E220000";
		ram_buffer(2207) := X"00000000";
		ram_buffer(2208) := X"10400018";
		ram_buffer(2209) := X"00101880";
		ram_buffer(2210) := X"00701021";
		ram_buffer(2211) := X"00021080";
		ram_buffer(2212) := X"02422021";
		ram_buffer(2213) := X"8C850004";
		ram_buffer(2214) := X"24420008";
		ram_buffer(2215) := X"8CA50004";
		ram_buffer(2216) := X"02421021";
		ram_buffer(2217) := X"14A20004";
		ram_buffer(2218) := X"AC850004";
		ram_buffer(2219) := X"8CA20004";
		ram_buffer(2220) := X"00000000";
		ram_buffer(2221) := X"AC820004";
		ram_buffer(2222) := X"00701821";
		ram_buffer(2223) := X"00031880";
		ram_buffer(2224) := X"02439021";
		ram_buffer(2225) := X"8E420004";
		ram_buffer(2226) := X"00000000";
		ram_buffer(2227) := X"8C42000C";
		ram_buffer(2228) := X"00000000";
		ram_buffer(2229) := X"AF82800C";
		ram_buffer(2230) := X"AF908030";
		ram_buffer(2231) := X"1000FFD5";
		ram_buffer(2232) := X"00000000";
		ram_buffer(2233) := X"16000003";
		ram_buffer(2234) := X"24050B05";
		ram_buffer(2235) := X"0C00023D";
		ram_buffer(2236) := X"02602025";
		ram_buffer(2237) := X"2610FFFF";
		ram_buffer(2238) := X"1000FFDF";
		ram_buffer(2239) := X"2631FFEC";
		ram_buffer(2240) := X"27BDFFE0";
		ram_buffer(2241) := X"AFB10018";
		ram_buffer(2242) := X"AFB00014";
		ram_buffer(2243) := X"AFBF001C";
		ram_buffer(2244) := X"00808025";
		ram_buffer(2245) := X"14800005";
		ram_buffer(2246) := X"00A08825";
		ram_buffer(2247) := X"3C040000";
		ram_buffer(2248) := X"24050B15";
		ram_buffer(2249) := X"0C00023D";
		ram_buffer(2250) := X"248445CC";
		ram_buffer(2251) := X"8F85800C";
		ram_buffer(2252) := X"02002025";
		ram_buffer(2253) := X"0C00026E";
		ram_buffer(2254) := X"24A50018";
		ram_buffer(2255) := X"8FBF001C";
		ram_buffer(2256) := X"8FB00014";
		ram_buffer(2257) := X"02202025";
		ram_buffer(2258) := X"8FB10018";
		ram_buffer(2259) := X"24050001";
		ram_buffer(2260) := X"0800075E";
		ram_buffer(2261) := X"27BD0020";
		ram_buffer(2262) := X"27BDFFE0";
		ram_buffer(2263) := X"AFB20018";
		ram_buffer(2264) := X"AFB10014";
		ram_buffer(2265) := X"AFB00010";
		ram_buffer(2266) := X"AFBF001C";
		ram_buffer(2267) := X"00808825";
		ram_buffer(2268) := X"00A08025";
		ram_buffer(2269) := X"14800005";
		ram_buffer(2270) := X"00C09025";
		ram_buffer(2271) := X"3C040000";
		ram_buffer(2272) := X"24050B26";
		ram_buffer(2273) := X"0C00023D";
		ram_buffer(2274) := X"248445CC";
		ram_buffer(2275) := X"8F828010";
		ram_buffer(2276) := X"00000000";
		ram_buffer(2277) := X"14400004";
		ram_buffer(2278) := X"3C040000";
		ram_buffer(2279) := X"24050B2A";
		ram_buffer(2280) := X"0C00023D";
		ram_buffer(2281) := X"248445CC";
		ram_buffer(2282) := X"8F82800C";
		ram_buffer(2283) := X"3C038000";
		ram_buffer(2284) := X"8F85800C";
		ram_buffer(2285) := X"02038025";
		ram_buffer(2286) := X"02202025";
		ram_buffer(2287) := X"AC500018";
		ram_buffer(2288) := X"0C000260";
		ram_buffer(2289) := X"24A50018";
		ram_buffer(2290) := X"8FBF001C";
		ram_buffer(2291) := X"8FB10014";
		ram_buffer(2292) := X"8FB00010";
		ram_buffer(2293) := X"02402025";
		ram_buffer(2294) := X"8FB20018";
		ram_buffer(2295) := X"24050001";
		ram_buffer(2296) := X"0800075E";
		ram_buffer(2297) := X"27BD0020";
		ram_buffer(2298) := X"8C82000C";
		ram_buffer(2299) := X"27BDFFE0";
		ram_buffer(2300) := X"AFB00014";
		ram_buffer(2301) := X"8C50000C";
		ram_buffer(2302) := X"AFBF001C";
		ram_buffer(2303) := X"16000005";
		ram_buffer(2304) := X"AFB10018";
		ram_buffer(2305) := X"3C040000";
		ram_buffer(2306) := X"24050B70";
		ram_buffer(2307) := X"0C00023D";
		ram_buffer(2308) := X"248445CC";
		ram_buffer(2309) := X"26110018";
		ram_buffer(2310) := X"0C000289";
		ram_buffer(2311) := X"02202025";
		ram_buffer(2312) := X"8F828010";
		ram_buffer(2313) := X"00000000";
		ram_buffer(2314) := X"14400022";
		ram_buffer(2315) := X"3C040000";
		ram_buffer(2316) := X"26110004";
		ram_buffer(2317) := X"0C000289";
		ram_buffer(2318) := X"02202025";
		ram_buffer(2319) := X"8E04002C";
		ram_buffer(2320) := X"8F828030";
		ram_buffer(2321) := X"00000000";
		ram_buffer(2322) := X"0044102B";
		ram_buffer(2323) := X"10400002";
		ram_buffer(2324) := X"00000000";
		ram_buffer(2325) := X"AF848030";
		ram_buffer(2326) := X"00041080";
		ram_buffer(2327) := X"00441021";
		ram_buffer(2328) := X"3C040000";
		ram_buffer(2329) := X"00021080";
		ram_buffer(2330) := X"248446E4";
		ram_buffer(2331) := X"02202825";
		ram_buffer(2332) := X"00822021";
		ram_buffer(2333) := X"0C000260";
		ram_buffer(2334) := X"00000000";
		ram_buffer(2335) := X"8F82800C";
		ram_buffer(2336) := X"8E03002C";
		ram_buffer(2337) := X"8C42002C";
		ram_buffer(2338) := X"00000000";
		ram_buffer(2339) := X"0043182B";
		ram_buffer(2340) := X"10600003";
		ram_buffer(2341) := X"00001025";
		ram_buffer(2342) := X"24020001";
		ram_buffer(2343) := X"AF828024";
		ram_buffer(2344) := X"8FBF001C";
		ram_buffer(2345) := X"8FB10018";
		ram_buffer(2346) := X"8FB00014";
		ram_buffer(2347) := X"03E00008";
		ram_buffer(2348) := X"27BD0020";
		ram_buffer(2349) := X"02202825";
		ram_buffer(2350) := X"1000FFEE";
		ram_buffer(2351) := X"248446A8";
		ram_buffer(2352) := X"8F828010";
		ram_buffer(2353) := X"27BDFFE0";
		ram_buffer(2354) := X"AFB10018";
		ram_buffer(2355) := X"AFB00014";
		ram_buffer(2356) := X"AFBF001C";
		ram_buffer(2357) := X"00808825";
		ram_buffer(2358) := X"14400005";
		ram_buffer(2359) := X"00A08025";
		ram_buffer(2360) := X"3C040000";
		ram_buffer(2361) := X"24050BA8";
		ram_buffer(2362) := X"0C00023D";
		ram_buffer(2363) := X"248445CC";
		ram_buffer(2364) := X"3C028000";
		ram_buffer(2365) := X"02028025";
		ram_buffer(2366) := X"AE300000";
		ram_buffer(2367) := X"8E30000C";
		ram_buffer(2368) := X"00000000";
		ram_buffer(2369) := X"16000004";
		ram_buffer(2370) := X"24050BB0";
		ram_buffer(2371) := X"3C040000";
		ram_buffer(2372) := X"0C00023D";
		ram_buffer(2373) := X"248445CC";
		ram_buffer(2374) := X"02202025";
		ram_buffer(2375) := X"0C000289";
		ram_buffer(2376) := X"26110004";
		ram_buffer(2377) := X"0C000289";
		ram_buffer(2378) := X"02202025";
		ram_buffer(2379) := X"8E04002C";
		ram_buffer(2380) := X"8F828030";
		ram_buffer(2381) := X"00000000";
		ram_buffer(2382) := X"0044102B";
		ram_buffer(2383) := X"10400002";
		ram_buffer(2384) := X"00000000";
		ram_buffer(2385) := X"AF848030";
		ram_buffer(2386) := X"00041080";
		ram_buffer(2387) := X"00441021";
		ram_buffer(2388) := X"3C040000";
		ram_buffer(2389) := X"00021080";
		ram_buffer(2390) := X"248446E4";
		ram_buffer(2391) := X"00822021";
		ram_buffer(2392) := X"0C000260";
		ram_buffer(2393) := X"02202825";
		ram_buffer(2394) := X"8F82800C";
		ram_buffer(2395) := X"8E03002C";
		ram_buffer(2396) := X"8C42002C";
		ram_buffer(2397) := X"00000000";
		ram_buffer(2398) := X"0043182B";
		ram_buffer(2399) := X"10600003";
		ram_buffer(2400) := X"00001025";
		ram_buffer(2401) := X"24020001";
		ram_buffer(2402) := X"AF828024";
		ram_buffer(2403) := X"8FBF001C";
		ram_buffer(2404) := X"8FB10018";
		ram_buffer(2405) := X"8FB00014";
		ram_buffer(2406) := X"03E00008";
		ram_buffer(2407) := X"27BD0020";
		ram_buffer(2408) := X"27BDFFE8";
		ram_buffer(2409) := X"AFB00010";
		ram_buffer(2410) := X"AFBF0014";
		ram_buffer(2411) := X"14800005";
		ram_buffer(2412) := X"00808025";
		ram_buffer(2413) := X"3C040000";
		ram_buffer(2414) := X"24050BD0";
		ram_buffer(2415) := X"0C00023D";
		ram_buffer(2416) := X"248445CC";
		ram_buffer(2417) := X"8F828020";
		ram_buffer(2418) := X"8FBF0014";
		ram_buffer(2419) := X"AE020000";
		ram_buffer(2420) := X"8F828034";
		ram_buffer(2421) := X"00000000";
		ram_buffer(2422) := X"AE020004";
		ram_buffer(2423) := X"8FB00010";
		ram_buffer(2424) := X"03E00008";
		ram_buffer(2425) := X"27BD0018";
		ram_buffer(2426) := X"24020001";
		ram_buffer(2427) := X"AF828024";
		ram_buffer(2428) := X"03E00008";
		ram_buffer(2429) := X"00000000";
		ram_buffer(2430) := X"14800003";
		ram_buffer(2431) := X"00000000";
		ram_buffer(2432) := X"8F84800C";
		ram_buffer(2433) := X"00000000";
		ram_buffer(2434) := X"8C840030";
		ram_buffer(2435) := X"240500A5";
		ram_buffer(2436) := X"00801825";
		ram_buffer(2437) := X"90660000";
		ram_buffer(2438) := X"00000000";
		ram_buffer(2439) := X"10C50004";
		ram_buffer(2440) := X"00641023";
		ram_buffer(2441) := X"00021082";
		ram_buffer(2442) := X"03E00008";
		ram_buffer(2443) := X"3042FFFF";
		ram_buffer(2444) := X"1000FFF8";
		ram_buffer(2445) := X"24630001";
		ram_buffer(2446) := X"8F82800C";
		ram_buffer(2447) := X"03E00008";
		ram_buffer(2448) := X"00000000";
		ram_buffer(2449) := X"8F83802C";
		ram_buffer(2450) := X"00000000";
		ram_buffer(2451) := X"10600005";
		ram_buffer(2452) := X"24020001";
		ram_buffer(2453) := X"8F828010";
		ram_buffer(2454) := X"00000000";
		ram_buffer(2455) := X"2C420001";
		ram_buffer(2456) := X"00021040";
		ram_buffer(2457) := X"03E00008";
		ram_buffer(2458) := X"00000000";
		ram_buffer(2459) := X"1080003E";
		ram_buffer(2460) := X"00000000";
		ram_buffer(2461) := X"8F82800C";
		ram_buffer(2462) := X"8C83002C";
		ram_buffer(2463) := X"8C42002C";
		ram_buffer(2464) := X"27BDFFE0";
		ram_buffer(2465) := X"0062102B";
		ram_buffer(2466) := X"AFBF001C";
		ram_buffer(2467) := X"AFB20018";
		ram_buffer(2468) := X"AFB10014";
		ram_buffer(2469) := X"1040002F";
		ram_buffer(2470) := X"AFB00010";
		ram_buffer(2471) := X"8C820018";
		ram_buffer(2472) := X"00000000";
		ram_buffer(2473) := X"04400008";
		ram_buffer(2474) := X"00031080";
		ram_buffer(2475) := X"8F82800C";
		ram_buffer(2476) := X"00000000";
		ram_buffer(2477) := X"8C45002C";
		ram_buffer(2478) := X"24020005";
		ram_buffer(2479) := X"00451023";
		ram_buffer(2480) := X"AC820018";
		ram_buffer(2481) := X"00031080";
		ram_buffer(2482) := X"00431021";
		ram_buffer(2483) := X"3C110000";
		ram_buffer(2484) := X"00021080";
		ram_buffer(2485) := X"263146E4";
		ram_buffer(2486) := X"8C830014";
		ram_buffer(2487) := X"02221021";
		ram_buffer(2488) := X"14620017";
		ram_buffer(2489) := X"24920004";
		ram_buffer(2490) := X"00808025";
		ram_buffer(2491) := X"0C000289";
		ram_buffer(2492) := X"02402025";
		ram_buffer(2493) := X"8F82800C";
		ram_buffer(2494) := X"8F838030";
		ram_buffer(2495) := X"8C42002C";
		ram_buffer(2496) := X"00000000";
		ram_buffer(2497) := X"0062182B";
		ram_buffer(2498) := X"10600002";
		ram_buffer(2499) := X"AE02002C";
		ram_buffer(2500) := X"AF828030";
		ram_buffer(2501) := X"00022080";
		ram_buffer(2502) := X"00822021";
		ram_buffer(2503) := X"00042080";
		ram_buffer(2504) := X"8FBF001C";
		ram_buffer(2505) := X"8FB00010";
		ram_buffer(2506) := X"02402825";
		ram_buffer(2507) := X"02242021";
		ram_buffer(2508) := X"8FB20018";
		ram_buffer(2509) := X"8FB10014";
		ram_buffer(2510) := X"08000260";
		ram_buffer(2511) := X"27BD0020";
		ram_buffer(2512) := X"8F82800C";
		ram_buffer(2513) := X"00000000";
		ram_buffer(2514) := X"8C42002C";
		ram_buffer(2515) := X"00000000";
		ram_buffer(2516) := X"AC82002C";
		ram_buffer(2517) := X"8FBF001C";
		ram_buffer(2518) := X"8FB20018";
		ram_buffer(2519) := X"8FB10014";
		ram_buffer(2520) := X"8FB00010";
		ram_buffer(2521) := X"27BD0020";
		ram_buffer(2522) := X"03E00008";
		ram_buffer(2523) := X"00000000";
		ram_buffer(2524) := X"14800009";
		ram_buffer(2525) := X"00001025";
		ram_buffer(2526) := X"03E00008";
		ram_buffer(2527) := X"00000000";
		ram_buffer(2528) := X"00001025";
		ram_buffer(2529) := X"8FBF001C";
		ram_buffer(2530) := X"8FB10018";
		ram_buffer(2531) := X"8FB00014";
		ram_buffer(2532) := X"03E00008";
		ram_buffer(2533) := X"27BD0020";
		ram_buffer(2534) := X"8F82800C";
		ram_buffer(2535) := X"27BDFFE0";
		ram_buffer(2536) := X"AFB00014";
		ram_buffer(2537) := X"AFBF001C";
		ram_buffer(2538) := X"AFB10018";
		ram_buffer(2539) := X"10820005";
		ram_buffer(2540) := X"00808025";
		ram_buffer(2541) := X"3C040000";
		ram_buffer(2542) := X"24050ED6";
		ram_buffer(2543) := X"0C00023D";
		ram_buffer(2544) := X"248445CC";
		ram_buffer(2545) := X"8E02004C";
		ram_buffer(2546) := X"00000000";
		ram_buffer(2547) := X"14400005";
		ram_buffer(2548) := X"3C040000";
		ram_buffer(2549) := X"24050ED8";
		ram_buffer(2550) := X"0C00023D";
		ram_buffer(2551) := X"248445CC";
		ram_buffer(2552) := X"8E02004C";
		ram_buffer(2553) := X"8E04002C";
		ram_buffer(2554) := X"8E030048";
		ram_buffer(2555) := X"2442FFFF";
		ram_buffer(2556) := X"1083FFE3";
		ram_buffer(2557) := X"AE02004C";
		ram_buffer(2558) := X"1440FFE2";
		ram_buffer(2559) := X"00001025";
		ram_buffer(2560) := X"26110004";
		ram_buffer(2561) := X"0C000289";
		ram_buffer(2562) := X"02202025";
		ram_buffer(2563) := X"8E040048";
		ram_buffer(2564) := X"24020005";
		ram_buffer(2565) := X"00441023";
		ram_buffer(2566) := X"AE020018";
		ram_buffer(2567) := X"8F828030";
		ram_buffer(2568) := X"00000000";
		ram_buffer(2569) := X"0044102B";
		ram_buffer(2570) := X"10400002";
		ram_buffer(2571) := X"AE04002C";
		ram_buffer(2572) := X"AF848030";
		ram_buffer(2573) := X"00041080";
		ram_buffer(2574) := X"00442021";
		ram_buffer(2575) := X"3C020000";
		ram_buffer(2576) := X"244246E4";
		ram_buffer(2577) := X"00042080";
		ram_buffer(2578) := X"00442021";
		ram_buffer(2579) := X"0C000260";
		ram_buffer(2580) := X"02202825";
		ram_buffer(2581) := X"1000FFCB";
		ram_buffer(2582) := X"24020001";
		ram_buffer(2583) := X"27BDFFE8";
		ram_buffer(2584) := X"AFBF0014";
		ram_buffer(2585) := X"0C000238";
		ram_buffer(2586) := X"00000000";
		ram_buffer(2587) := X"8F82802C";
		ram_buffer(2588) := X"00000000";
		ram_buffer(2589) := X"10400008";
		ram_buffer(2590) := X"00000000";
		ram_buffer(2591) := X"8F83800C";
		ram_buffer(2592) := X"00000000";
		ram_buffer(2593) := X"8C620044";
		ram_buffer(2594) := X"00000000";
		ram_buffer(2595) := X"24420001";
		ram_buffer(2596) := X"AC620044";
		ram_buffer(2597) := X"8F82800C";
		ram_buffer(2598) := X"8FBF0014";
		ram_buffer(2599) := X"00000000";
		ram_buffer(2600) := X"03E00008";
		ram_buffer(2601) := X"27BD0018";
		ram_buffer(2602) := X"8F82802C";
		ram_buffer(2603) := X"00000000";
		ram_buffer(2604) := X"10400015";
		ram_buffer(2605) := X"00000000";
		ram_buffer(2606) := X"8F82800C";
		ram_buffer(2607) := X"00000000";
		ram_buffer(2608) := X"8C420044";
		ram_buffer(2609) := X"00000000";
		ram_buffer(2610) := X"1040000F";
		ram_buffer(2611) := X"00000000";
		ram_buffer(2612) := X"8F83800C";
		ram_buffer(2613) := X"00000000";
		ram_buffer(2614) := X"8C620044";
		ram_buffer(2615) := X"00000000";
		ram_buffer(2616) := X"2442FFFF";
		ram_buffer(2617) := X"AC620044";
		ram_buffer(2618) := X"8F82800C";
		ram_buffer(2619) := X"00000000";
		ram_buffer(2620) := X"8C420044";
		ram_buffer(2621) := X"00000000";
		ram_buffer(2622) := X"14400003";
		ram_buffer(2623) := X"00000000";
		ram_buffer(2624) := X"08000233";
		ram_buffer(2625) := X"00000000";
		ram_buffer(2626) := X"03E00008";
		ram_buffer(2627) := X"00000000";
		ram_buffer(2628) := X"27BDFFC8";
		ram_buffer(2629) := X"AFB2001C";
		ram_buffer(2630) := X"00069080";
		ram_buffer(2631) := X"AFB40024";
		ram_buffer(2632) := X"0080A025";
		ram_buffer(2633) := X"02402025";
		ram_buffer(2634) := X"AFB70030";
		ram_buffer(2635) := X"AFB50028";
		ram_buffer(2636) := X"AFB30020";
		ram_buffer(2637) := X"AFB10018";
		ram_buffer(2638) := X"AFBF0034";
		ram_buffer(2639) := X"AFB6002C";
		ram_buffer(2640) := X"AFB00014";
		ram_buffer(2641) := X"00A08825";
		ram_buffer(2642) := X"8FB3004C";
		ram_buffer(2643) := X"0C001008";
		ram_buffer(2644) := X"00E0A825";
		ram_buffer(2645) := X"1040008F";
		ram_buffer(2646) := X"2417FFFF";
		ram_buffer(2647) := X"24040058";
		ram_buffer(2648) := X"0C001008";
		ram_buffer(2649) := X"0040B025";
		ram_buffer(2650) := X"10400087";
		ram_buffer(2651) := X"00408025";
		ram_buffer(2652) := X"02403025";
		ram_buffer(2653) := X"240500A5";
		ram_buffer(2654) := X"AC560030";
		ram_buffer(2655) := X"0C001119";
		ram_buffer(2656) := X"02C02025";
		ram_buffer(2657) := X"2642FFFC";
		ram_buffer(2658) := X"8E120030";
		ram_buffer(2659) := X"02202825";
		ram_buffer(2660) := X"02429021";
		ram_buffer(2661) := X"2402FFFC";
		ram_buffer(2662) := X"02429024";
		ram_buffer(2663) := X"26230010";
		ram_buffer(2664) := X"26020034";
		ram_buffer(2665) := X"80A40000";
		ram_buffer(2666) := X"00000000";
		ram_buffer(2667) := X"A0440000";
		ram_buffer(2668) := X"80A40000";
		ram_buffer(2669) := X"00000000";
		ram_buffer(2670) := X"10800003";
		ram_buffer(2671) := X"24A50001";
		ram_buffer(2672) := X"1465FFF8";
		ram_buffer(2673) := X"24420001";
		ram_buffer(2674) := X"8FB60048";
		ram_buffer(2675) := X"00000000";
		ram_buffer(2676) := X"2EC20005";
		ram_buffer(2677) := X"14400002";
		ram_buffer(2678) := X"A2000043";
		ram_buffer(2679) := X"24160004";
		ram_buffer(2680) := X"26110004";
		ram_buffer(2681) := X"AE16002C";
		ram_buffer(2682) := X"AE160048";
		ram_buffer(2683) := X"02202025";
		ram_buffer(2684) := X"0C00025E";
		ram_buffer(2685) := X"AE00004C";
		ram_buffer(2686) := X"0C00025E";
		ram_buffer(2687) := X"26040018";
		ram_buffer(2688) := X"24020005";
		ram_buffer(2689) := X"0056B023";
		ram_buffer(2690) := X"AE000050";
		ram_buffer(2691) := X"AE100010";
		ram_buffer(2692) := X"AE160018";
		ram_buffer(2693) := X"AE100024";
		ram_buffer(2694) := X"AE000044";
		ram_buffer(2695) := X"A2000054";
		ram_buffer(2696) := X"A2000055";
		ram_buffer(2697) := X"02A03025";
		ram_buffer(2698) := X"02802825";
		ram_buffer(2699) := X"0C0000FA";
		ram_buffer(2700) := X"02402025";
		ram_buffer(2701) := X"12600002";
		ram_buffer(2702) := X"AE020000";
		ram_buffer(2703) := X"AE700000";
		ram_buffer(2704) := X"0C000A17";
		ram_buffer(2705) := X"00000000";
		ram_buffer(2706) := X"8F828038";
		ram_buffer(2707) := X"3C120000";
		ram_buffer(2708) := X"24420001";
		ram_buffer(2709) := X"AF828038";
		ram_buffer(2710) := X"8F82800C";
		ram_buffer(2711) := X"00000000";
		ram_buffer(2712) := X"14400058";
		ram_buffer(2713) := X"00000000";
		ram_buffer(2714) := X"AF90800C";
		ram_buffer(2715) := X"8F838038";
		ram_buffer(2716) := X"24020001";
		ram_buffer(2717) := X"14620022";
		ram_buffer(2718) := X"00000000";
		ram_buffer(2719) := X"0C000256";
		ram_buffer(2720) := X"264446E4";
		ram_buffer(2721) := X"3C040000";
		ram_buffer(2722) := X"0C000256";
		ram_buffer(2723) := X"248446F8";
		ram_buffer(2724) := X"3C040000";
		ram_buffer(2725) := X"0C000256";
		ram_buffer(2726) := X"2484470C";
		ram_buffer(2727) := X"3C040000";
		ram_buffer(2728) := X"0C000256";
		ram_buffer(2729) := X"24844720";
		ram_buffer(2730) := X"3C040000";
		ram_buffer(2731) := X"24844734";
		ram_buffer(2732) := X"0C000256";
		ram_buffer(2733) := X"3C140000";
		ram_buffer(2734) := X"3C130000";
		ram_buffer(2735) := X"0C000256";
		ram_buffer(2736) := X"268446D0";
		ram_buffer(2737) := X"0C000256";
		ram_buffer(2738) := X"266446BC";
		ram_buffer(2739) := X"3C040000";
		ram_buffer(2740) := X"0C000256";
		ram_buffer(2741) := X"248446A8";
		ram_buffer(2742) := X"3C040000";
		ram_buffer(2743) := X"0C000256";
		ram_buffer(2744) := X"24844694";
		ram_buffer(2745) := X"3C040000";
		ram_buffer(2746) := X"24844680";
		ram_buffer(2747) := X"269446D0";
		ram_buffer(2748) := X"0C000256";
		ram_buffer(2749) := X"267346BC";
		ram_buffer(2750) := X"AF948044";
		ram_buffer(2751) := X"AF938040";
		ram_buffer(2752) := X"8F82801C";
		ram_buffer(2753) := X"8E04002C";
		ram_buffer(2754) := X"24420001";
		ram_buffer(2755) := X"AF82801C";
		ram_buffer(2756) := X"8F828030";
		ram_buffer(2757) := X"00000000";
		ram_buffer(2758) := X"0044102B";
		ram_buffer(2759) := X"10400003";
		ram_buffer(2760) := X"00041080";
		ram_buffer(2761) := X"AF848030";
		ram_buffer(2762) := X"00041080";
		ram_buffer(2763) := X"00441021";
		ram_buffer(2764) := X"00021080";
		ram_buffer(2765) := X"264446E4";
		ram_buffer(2766) := X"00822021";
		ram_buffer(2767) := X"0C000260";
		ram_buffer(2768) := X"02202825";
		ram_buffer(2769) := X"0C000A2A";
		ram_buffer(2770) := X"00000000";
		ram_buffer(2771) := X"8F82802C";
		ram_buffer(2772) := X"00000000";
		ram_buffer(2773) := X"1040000F";
		ram_buffer(2774) := X"24170001";
		ram_buffer(2775) := X"8F82800C";
		ram_buffer(2776) := X"8E03002C";
		ram_buffer(2777) := X"8C42002C";
		ram_buffer(2778) := X"00000000";
		ram_buffer(2779) := X"0043102B";
		ram_buffer(2780) := X"10400008";
		ram_buffer(2781) := X"00000000";
		ram_buffer(2782) := X"0C00017D";
		ram_buffer(2783) := X"00000000";
		ram_buffer(2784) := X"10000004";
		ram_buffer(2785) := X"00000000";
		ram_buffer(2786) := X"0C001030";
		ram_buffer(2787) := X"02C02025";
		ram_buffer(2788) := X"2417FFFF";
		ram_buffer(2789) := X"8FBF0034";
		ram_buffer(2790) := X"02E01025";
		ram_buffer(2791) := X"8FB6002C";
		ram_buffer(2792) := X"8FB70030";
		ram_buffer(2793) := X"8FB50028";
		ram_buffer(2794) := X"8FB40024";
		ram_buffer(2795) := X"8FB30020";
		ram_buffer(2796) := X"8FB2001C";
		ram_buffer(2797) := X"8FB10018";
		ram_buffer(2798) := X"8FB00014";
		ram_buffer(2799) := X"03E00008";
		ram_buffer(2800) := X"27BD0038";
		ram_buffer(2801) := X"8F82802C";
		ram_buffer(2802) := X"00000000";
		ram_buffer(2803) := X"1440FFCC";
		ram_buffer(2804) := X"00000000";
		ram_buffer(2805) := X"8F82800C";
		ram_buffer(2806) := X"8E03002C";
		ram_buffer(2807) := X"8C42002C";
		ram_buffer(2808) := X"00000000";
		ram_buffer(2809) := X"0062102B";
		ram_buffer(2810) := X"1440FFC5";
		ram_buffer(2811) := X"00000000";
		ram_buffer(2812) := X"AF90800C";
		ram_buffer(2813) := X"1000FFC2";
		ram_buffer(2814) := X"00000000";
		ram_buffer(2815) := X"27BDFFE0";
		ram_buffer(2816) := X"27828014";
		ram_buffer(2817) := X"3C050000";
		ram_buffer(2818) := X"3C040000";
		ram_buffer(2819) := X"00003825";
		ram_buffer(2820) := X"AFA20014";
		ram_buffer(2821) := X"AFA00010";
		ram_buffer(2822) := X"2406012C";
		ram_buffer(2823) := X"24A545E4";
		ram_buffer(2824) := X"AFB00018";
		ram_buffer(2825) := X"AFBF001C";
		ram_buffer(2826) := X"0C000A44";
		ram_buffer(2827) := X"248435F4";
		ram_buffer(2828) := X"00408025";
		ram_buffer(2829) := X"24020001";
		ram_buffer(2830) := X"1602000C";
		ram_buffer(2831) := X"2402FFFF";
		ram_buffer(2832) := X"0C000238";
		ram_buffer(2833) := X"00000000";
		ram_buffer(2834) := X"2402FFFF";
		ram_buffer(2835) := X"AF828018";
		ram_buffer(2836) := X"8FBF001C";
		ram_buffer(2837) := X"AF90802C";
		ram_buffer(2838) := X"8FB00018";
		ram_buffer(2839) := X"27BD0020";
		ram_buffer(2840) := X"AF808034";
		ram_buffer(2841) := X"08000FF8";
		ram_buffer(2842) := X"00000000";
		ram_buffer(2843) := X"16020007";
		ram_buffer(2844) := X"3C040000";
		ram_buffer(2845) := X"8FBF001C";
		ram_buffer(2846) := X"8FB00018";
		ram_buffer(2847) := X"2405078B";
		ram_buffer(2848) := X"248445CC";
		ram_buffer(2849) := X"0800023D";
		ram_buffer(2850) := X"27BD0020";
		ram_buffer(2851) := X"8FBF001C";
		ram_buffer(2852) := X"8FB00018";
		ram_buffer(2853) := X"03E00008";
		ram_buffer(2854) := X"27BD0020";
		ram_buffer(2855) := X"27BDFFE0";
		ram_buffer(2856) := X"AFB00014";
		ram_buffer(2857) := X"00808025";
		ram_buffer(2858) := X"AFBF001C";
		ram_buffer(2859) := X"0C000A17";
		ram_buffer(2860) := X"AFB10018";
		ram_buffer(2861) := X"16000004";
		ram_buffer(2862) := X"26110004";
		ram_buffer(2863) := X"8F90800C";
		ram_buffer(2864) := X"00000000";
		ram_buffer(2865) := X"26110004";
		ram_buffer(2866) := X"0C000289";
		ram_buffer(2867) := X"02202025";
		ram_buffer(2868) := X"8E020028";
		ram_buffer(2869) := X"00000000";
		ram_buffer(2870) := X"10400003";
		ram_buffer(2871) := X"00000000";
		ram_buffer(2872) := X"0C000289";
		ram_buffer(2873) := X"26040018";
		ram_buffer(2874) := X"8F82801C";
		ram_buffer(2875) := X"00000000";
		ram_buffer(2876) := X"24420001";
		ram_buffer(2877) := X"AF82801C";
		ram_buffer(2878) := X"8F82800C";
		ram_buffer(2879) := X"00000000";
		ram_buffer(2880) := X"1602001E";
		ram_buffer(2881) := X"02202825";
		ram_buffer(2882) := X"3C040000";
		ram_buffer(2883) := X"0C000260";
		ram_buffer(2884) := X"24844694";
		ram_buffer(2885) := X"8F82803C";
		ram_buffer(2886) := X"00000000";
		ram_buffer(2887) := X"24420001";
		ram_buffer(2888) := X"AF82803C";
		ram_buffer(2889) := X"0C000A2A";
		ram_buffer(2890) := X"00000000";
		ram_buffer(2891) := X"8F82802C";
		ram_buffer(2892) := X"00000000";
		ram_buffer(2893) := X"1040001D";
		ram_buffer(2894) := X"00000000";
		ram_buffer(2895) := X"8F82800C";
		ram_buffer(2896) := X"00000000";
		ram_buffer(2897) := X"16020019";
		ram_buffer(2898) := X"00000000";
		ram_buffer(2899) := X"8F828010";
		ram_buffer(2900) := X"00000000";
		ram_buffer(2901) := X"10400004";
		ram_buffer(2902) := X"24050465";
		ram_buffer(2903) := X"3C040000";
		ram_buffer(2904) := X"0C00023D";
		ram_buffer(2905) := X"248445CC";
		ram_buffer(2906) := X"8FBF001C";
		ram_buffer(2907) := X"8FB10018";
		ram_buffer(2908) := X"8FB00014";
		ram_buffer(2909) := X"0800017D";
		ram_buffer(2910) := X"27BD0020";
		ram_buffer(2911) := X"8F828038";
		ram_buffer(2912) := X"8E040030";
		ram_buffer(2913) := X"2442FFFF";
		ram_buffer(2914) := X"AF828038";
		ram_buffer(2915) := X"0C001030";
		ram_buffer(2916) := X"00000000";
		ram_buffer(2917) := X"0C001030";
		ram_buffer(2918) := X"02002025";
		ram_buffer(2919) := X"0C000733";
		ram_buffer(2920) := X"00000000";
		ram_buffer(2921) := X"1000FFDF";
		ram_buffer(2922) := X"00000000";
		ram_buffer(2923) := X"8FBF001C";
		ram_buffer(2924) := X"8FB10018";
		ram_buffer(2925) := X"8FB00014";
		ram_buffer(2926) := X"03E00008";
		ram_buffer(2927) := X"27BD0020";
		ram_buffer(2928) := X"27BDFFE0";
		ram_buffer(2929) := X"AFB10018";
		ram_buffer(2930) := X"AFBF001C";
		ram_buffer(2931) := X"AFB00014";
		ram_buffer(2932) := X"14800005";
		ram_buffer(2933) := X"00808825";
		ram_buffer(2934) := X"3C040000";
		ram_buffer(2935) := X"24050502";
		ram_buffer(2936) := X"0C00023D";
		ram_buffer(2937) := X"248445CC";
		ram_buffer(2938) := X"8F83800C";
		ram_buffer(2939) := X"00000000";
		ram_buffer(2940) := X"12230016";
		ram_buffer(2941) := X"00001025";
		ram_buffer(2942) := X"0C000A17";
		ram_buffer(2943) := X"00000000";
		ram_buffer(2944) := X"8E300014";
		ram_buffer(2945) := X"0C000A2A";
		ram_buffer(2946) := X"00000000";
		ram_buffer(2947) := X"8F838044";
		ram_buffer(2948) := X"00000000";
		ram_buffer(2949) := X"1203000D";
		ram_buffer(2950) := X"24020002";
		ram_buffer(2951) := X"8F838040";
		ram_buffer(2952) := X"00000000";
		ram_buffer(2953) := X"12030009";
		ram_buffer(2954) := X"00000000";
		ram_buffer(2955) := X"3C020000";
		ram_buffer(2956) := X"24424680";
		ram_buffer(2957) := X"1602000A";
		ram_buffer(2958) := X"3C030000";
		ram_buffer(2959) := X"8E220028";
		ram_buffer(2960) := X"00000000";
		ram_buffer(2961) := X"2C420001";
		ram_buffer(2962) := X"24420002";
		ram_buffer(2963) := X"8FBF001C";
		ram_buffer(2964) := X"8FB10018";
		ram_buffer(2965) := X"8FB00014";
		ram_buffer(2966) := X"03E00008";
		ram_buffer(2967) := X"27BD0020";
		ram_buffer(2968) := X"24634694";
		ram_buffer(2969) := X"1203FFF9";
		ram_buffer(2970) := X"24020004";
		ram_buffer(2971) := X"1200FFF7";
		ram_buffer(2972) := X"00000000";
		ram_buffer(2973) := X"1000FFF5";
		ram_buffer(2974) := X"24020001";
		ram_buffer(2975) := X"27BDFFE8";
		ram_buffer(2976) := X"AFB00010";
		ram_buffer(2977) := X"AFBF0014";
		ram_buffer(2978) := X"0C000A17";
		ram_buffer(2979) := X"00808025";
		ram_buffer(2980) := X"16000003";
		ram_buffer(2981) := X"02002025";
		ram_buffer(2982) := X"8F84800C";
		ram_buffer(2983) := X"00000000";
		ram_buffer(2984) := X"8C90002C";
		ram_buffer(2985) := X"0C000A2A";
		ram_buffer(2986) := X"00000000";
		ram_buffer(2987) := X"8FBF0014";
		ram_buffer(2988) := X"02001025";
		ram_buffer(2989) := X"8FB00010";
		ram_buffer(2990) := X"03E00008";
		ram_buffer(2991) := X"27BD0018";
		ram_buffer(2992) := X"27BDFFD8";
		ram_buffer(2993) := X"2CA20005";
		ram_buffer(2994) := X"AFB2001C";
		ram_buffer(2995) := X"AFB00014";
		ram_buffer(2996) := X"AFBF0024";
		ram_buffer(2997) := X"AFB30020";
		ram_buffer(2998) := X"AFB10018";
		ram_buffer(2999) := X"00808025";
		ram_buffer(3000) := X"14400006";
		ram_buffer(3001) := X"00A09025";
		ram_buffer(3002) := X"3C040000";
		ram_buffer(3003) := X"24050587";
		ram_buffer(3004) := X"0C00023D";
		ram_buffer(3005) := X"248445CC";
		ram_buffer(3006) := X"24120004";
		ram_buffer(3007) := X"0C000A17";
		ram_buffer(3008) := X"00000000";
		ram_buffer(3009) := X"16000003";
		ram_buffer(3010) := X"00000000";
		ram_buffer(3011) := X"8F90800C";
		ram_buffer(3012) := X"00000000";
		ram_buffer(3013) := X"8E020048";
		ram_buffer(3014) := X"00000000";
		ram_buffer(3015) := X"12420035";
		ram_buffer(3016) := X"0052182B";
		ram_buffer(3017) := X"1060003A";
		ram_buffer(3018) := X"00000000";
		ram_buffer(3019) := X"8F83800C";
		ram_buffer(3020) := X"00000000";
		ram_buffer(3021) := X"12030007";
		ram_buffer(3022) := X"00008825";
		ram_buffer(3023) := X"8F83800C";
		ram_buffer(3024) := X"00000000";
		ram_buffer(3025) := X"8C71002C";
		ram_buffer(3026) := X"00000000";
		ram_buffer(3027) := X"0251882B";
		ram_buffer(3028) := X"3A310001";
		ram_buffer(3029) := X"8E03002C";
		ram_buffer(3030) := X"00000000";
		ram_buffer(3031) := X"14430002";
		ram_buffer(3032) := X"00000000";
		ram_buffer(3033) := X"AE12002C";
		ram_buffer(3034) := X"8E020018";
		ram_buffer(3035) := X"00000000";
		ram_buffer(3036) := X"04400004";
		ram_buffer(3037) := X"AE120048";
		ram_buffer(3038) := X"24050005";
		ram_buffer(3039) := X"00B29023";
		ram_buffer(3040) := X"AE120018";
		ram_buffer(3041) := X"00031080";
		ram_buffer(3042) := X"00431021";
		ram_buffer(3043) := X"3C120000";
		ram_buffer(3044) := X"00021080";
		ram_buffer(3045) := X"265246E4";
		ram_buffer(3046) := X"8E030014";
		ram_buffer(3047) := X"02421021";
		ram_buffer(3048) := X"14620010";
		ram_buffer(3049) := X"26130004";
		ram_buffer(3050) := X"0C000289";
		ram_buffer(3051) := X"02602025";
		ram_buffer(3052) := X"8E02002C";
		ram_buffer(3053) := X"8F838030";
		ram_buffer(3054) := X"00000000";
		ram_buffer(3055) := X"0062182B";
		ram_buffer(3056) := X"10600002";
		ram_buffer(3057) := X"00000000";
		ram_buffer(3058) := X"AF828030";
		ram_buffer(3059) := X"00022080";
		ram_buffer(3060) := X"00822021";
		ram_buffer(3061) := X"00042080";
		ram_buffer(3062) := X"02602825";
		ram_buffer(3063) := X"0C000260";
		ram_buffer(3064) := X"02442021";
		ram_buffer(3065) := X"12200003";
		ram_buffer(3066) := X"00000000";
		ram_buffer(3067) := X"0C00017D";
		ram_buffer(3068) := X"00000000";
		ram_buffer(3069) := X"8FBF0024";
		ram_buffer(3070) := X"8FB30020";
		ram_buffer(3071) := X"8FB2001C";
		ram_buffer(3072) := X"8FB10018";
		ram_buffer(3073) := X"8FB00014";
		ram_buffer(3074) := X"08000A2A";
		ram_buffer(3075) := X"27BD0028";
		ram_buffer(3076) := X"8F91800C";
		ram_buffer(3077) := X"00000000";
		ram_buffer(3078) := X"02118826";
		ram_buffer(3079) := X"1000FFCD";
		ram_buffer(3080) := X"2E310001";
		ram_buffer(3081) := X"27BDFFE0";
		ram_buffer(3082) := X"AFB00014";
		ram_buffer(3083) := X"00808025";
		ram_buffer(3084) := X"AFBF001C";
		ram_buffer(3085) := X"0C000A17";
		ram_buffer(3086) := X"AFB10018";
		ram_buffer(3087) := X"16000004";
		ram_buffer(3088) := X"26110004";
		ram_buffer(3089) := X"8F90800C";
		ram_buffer(3090) := X"00000000";
		ram_buffer(3091) := X"26110004";
		ram_buffer(3092) := X"0C000289";
		ram_buffer(3093) := X"02202025";
		ram_buffer(3094) := X"8E020028";
		ram_buffer(3095) := X"00000000";
		ram_buffer(3096) := X"10400004";
		ram_buffer(3097) := X"02202825";
		ram_buffer(3098) := X"0C000289";
		ram_buffer(3099) := X"26040018";
		ram_buffer(3100) := X"02202825";
		ram_buffer(3101) := X"3C110000";
		ram_buffer(3102) := X"0C000260";
		ram_buffer(3103) := X"26244680";
		ram_buffer(3104) := X"0C000A2A";
		ram_buffer(3105) := X"00000000";
		ram_buffer(3106) := X"8F82802C";
		ram_buffer(3107) := X"00000000";
		ram_buffer(3108) := X"10400007";
		ram_buffer(3109) := X"00000000";
		ram_buffer(3110) := X"0C000A17";
		ram_buffer(3111) := X"00000000";
		ram_buffer(3112) := X"0C000733";
		ram_buffer(3113) := X"00000000";
		ram_buffer(3114) := X"0C000A2A";
		ram_buffer(3115) := X"00000000";
		ram_buffer(3116) := X"8F82800C";
		ram_buffer(3117) := X"00000000";
		ram_buffer(3118) := X"16020017";
		ram_buffer(3119) := X"00000000";
		ram_buffer(3120) := X"8F82802C";
		ram_buffer(3121) := X"00000000";
		ram_buffer(3122) := X"1040000D";
		ram_buffer(3123) := X"00000000";
		ram_buffer(3124) := X"8F828010";
		ram_buffer(3125) := X"00000000";
		ram_buffer(3126) := X"10400004";
		ram_buffer(3127) := X"3C040000";
		ram_buffer(3128) := X"2405065E";
		ram_buffer(3129) := X"0C00023D";
		ram_buffer(3130) := X"248445CC";
		ram_buffer(3131) := X"8FBF001C";
		ram_buffer(3132) := X"8FB10018";
		ram_buffer(3133) := X"8FB00014";
		ram_buffer(3134) := X"0800017D";
		ram_buffer(3135) := X"27BD0020";
		ram_buffer(3136) := X"8F828038";
		ram_buffer(3137) := X"8E234680";
		ram_buffer(3138) := X"00000000";
		ram_buffer(3139) := X"14620007";
		ram_buffer(3140) := X"00000000";
		ram_buffer(3141) := X"AF80800C";
		ram_buffer(3142) := X"8FBF001C";
		ram_buffer(3143) := X"8FB10018";
		ram_buffer(3144) := X"8FB00014";
		ram_buffer(3145) := X"03E00008";
		ram_buffer(3146) := X"27BD0020";
		ram_buffer(3147) := X"8FBF001C";
		ram_buffer(3148) := X"8FB10018";
		ram_buffer(3149) := X"8FB00014";
		ram_buffer(3150) := X"08000883";
		ram_buffer(3151) := X"27BD0020";
		ram_buffer(3152) := X"14800029";
		ram_buffer(3153) := X"240506B2";
		ram_buffer(3154) := X"3C040000";
		ram_buffer(3155) := X"0800023D";
		ram_buffer(3156) := X"248445CC";
		ram_buffer(3157) := X"0C000A17";
		ram_buffer(3158) := X"00808025";
		ram_buffer(3159) := X"0C000746";
		ram_buffer(3160) := X"02002025";
		ram_buffer(3161) := X"1040001B";
		ram_buffer(3162) := X"26110004";
		ram_buffer(3163) := X"0C000289";
		ram_buffer(3164) := X"02202025";
		ram_buffer(3165) := X"8E04002C";
		ram_buffer(3166) := X"8F828030";
		ram_buffer(3167) := X"00000000";
		ram_buffer(3168) := X"0044102B";
		ram_buffer(3169) := X"10400003";
		ram_buffer(3170) := X"00041080";
		ram_buffer(3171) := X"AF848030";
		ram_buffer(3172) := X"00041080";
		ram_buffer(3173) := X"00441021";
		ram_buffer(3174) := X"3C040000";
		ram_buffer(3175) := X"00021080";
		ram_buffer(3176) := X"248446E4";
		ram_buffer(3177) := X"00822021";
		ram_buffer(3178) := X"0C000260";
		ram_buffer(3179) := X"02202825";
		ram_buffer(3180) := X"8F83800C";
		ram_buffer(3181) := X"8E02002C";
		ram_buffer(3182) := X"8C63002C";
		ram_buffer(3183) := X"00000000";
		ram_buffer(3184) := X"0043102B";
		ram_buffer(3185) := X"14400003";
		ram_buffer(3186) := X"00000000";
		ram_buffer(3187) := X"0C00017D";
		ram_buffer(3188) := X"00000000";
		ram_buffer(3189) := X"8FBF001C";
		ram_buffer(3190) := X"8FB10018";
		ram_buffer(3191) := X"8FB00014";
		ram_buffer(3192) := X"08000A2A";
		ram_buffer(3193) := X"27BD0020";
		ram_buffer(3194) := X"8F82800C";
		ram_buffer(3195) := X"27BDFFE0";
		ram_buffer(3196) := X"AFBF001C";
		ram_buffer(3197) := X"AFB10018";
		ram_buffer(3198) := X"1482FFD6";
		ram_buffer(3199) := X"AFB00014";
		ram_buffer(3200) := X"8FBF001C";
		ram_buffer(3201) := X"8FB10018";
		ram_buffer(3202) := X"8FB00014";
		ram_buffer(3203) := X"03E00008";
		ram_buffer(3204) := X"27BD0020";
		ram_buffer(3205) := X"8F828010";
		ram_buffer(3206) := X"27BDFFD0";
		ram_buffer(3207) := X"AFBF002C";
		ram_buffer(3208) := X"AFB50028";
		ram_buffer(3209) := X"AFB40024";
		ram_buffer(3210) := X"AFB30020";
		ram_buffer(3211) := X"AFB2001C";
		ram_buffer(3212) := X"AFB10018";
		ram_buffer(3213) := X"14400005";
		ram_buffer(3214) := X"AFB00014";
		ram_buffer(3215) := X"3C040000";
		ram_buffer(3216) := X"240507EF";
		ram_buffer(3217) := X"0C00023D";
		ram_buffer(3218) := X"248445CC";
		ram_buffer(3219) := X"0C000A17";
		ram_buffer(3220) := X"00000000";
		ram_buffer(3221) := X"8F828010";
		ram_buffer(3222) := X"00000000";
		ram_buffer(3223) := X"2442FFFF";
		ram_buffer(3224) := X"AF828010";
		ram_buffer(3225) := X"8F828010";
		ram_buffer(3226) := X"00000000";
		ram_buffer(3227) := X"1040000E";
		ram_buffer(3228) := X"00000000";
		ram_buffer(3229) := X"00008025";
		ram_buffer(3230) := X"0C000A2A";
		ram_buffer(3231) := X"00000000";
		ram_buffer(3232) := X"8FBF002C";
		ram_buffer(3233) := X"02001025";
		ram_buffer(3234) := X"8FB50028";
		ram_buffer(3235) := X"8FB40024";
		ram_buffer(3236) := X"8FB30020";
		ram_buffer(3237) := X"8FB2001C";
		ram_buffer(3238) := X"8FB10018";
		ram_buffer(3239) := X"8FB00014";
		ram_buffer(3240) := X"03E00008";
		ram_buffer(3241) := X"27BD0030";
		ram_buffer(3242) := X"8F828038";
		ram_buffer(3243) := X"00000000";
		ram_buffer(3244) := X"1040FFF0";
		ram_buffer(3245) := X"3C140000";
		ram_buffer(3246) := X"3C110000";
		ram_buffer(3247) := X"00008025";
		ram_buffer(3248) := X"269246A8";
		ram_buffer(3249) := X"263146E4";
		ram_buffer(3250) := X"24130001";
		ram_buffer(3251) := X"8E8246A8";
		ram_buffer(3252) := X"00000000";
		ram_buffer(3253) := X"1440001A";
		ram_buffer(3254) := X"00000000";
		ram_buffer(3255) := X"12000003";
		ram_buffer(3256) := X"00000000";
		ram_buffer(3257) := X"0C000733";
		ram_buffer(3258) := X"00000000";
		ram_buffer(3259) := X"8F908028";
		ram_buffer(3260) := X"00000000";
		ram_buffer(3261) := X"1200000A";
		ram_buffer(3262) := X"24110001";
		ram_buffer(3263) := X"0C000808";
		ram_buffer(3264) := X"00000000";
		ram_buffer(3265) := X"10400002";
		ram_buffer(3266) := X"00000000";
		ram_buffer(3267) := X"AF918024";
		ram_buffer(3268) := X"2610FFFF";
		ram_buffer(3269) := X"1600FFF9";
		ram_buffer(3270) := X"00000000";
		ram_buffer(3271) := X"AF808028";
		ram_buffer(3272) := X"8F828024";
		ram_buffer(3273) := X"00000000";
		ram_buffer(3274) := X"1040FFD2";
		ram_buffer(3275) := X"00000000";
		ram_buffer(3276) := X"0C00017D";
		ram_buffer(3277) := X"24100001";
		ram_buffer(3278) := X"1000FFCF";
		ram_buffer(3279) := X"00000000";
		ram_buffer(3280) := X"8E42000C";
		ram_buffer(3281) := X"00000000";
		ram_buffer(3282) := X"8C50000C";
		ram_buffer(3283) := X"00000000";
		ram_buffer(3284) := X"26040018";
		ram_buffer(3285) := X"0C000289";
		ram_buffer(3286) := X"26150004";
		ram_buffer(3287) := X"0C000289";
		ram_buffer(3288) := X"02A02025";
		ram_buffer(3289) := X"8E02002C";
		ram_buffer(3290) := X"8F838030";
		ram_buffer(3291) := X"00000000";
		ram_buffer(3292) := X"0062182B";
		ram_buffer(3293) := X"10600002";
		ram_buffer(3294) := X"00000000";
		ram_buffer(3295) := X"AF828030";
		ram_buffer(3296) := X"00022080";
		ram_buffer(3297) := X"00822021";
		ram_buffer(3298) := X"00042080";
		ram_buffer(3299) := X"02A02825";
		ram_buffer(3300) := X"0C000260";
		ram_buffer(3301) := X"02242021";
		ram_buffer(3302) := X"8F83800C";
		ram_buffer(3303) := X"8E02002C";
		ram_buffer(3304) := X"8C63002C";
		ram_buffer(3305) := X"00000000";
		ram_buffer(3306) := X"0043102B";
		ram_buffer(3307) := X"1440FFC7";
		ram_buffer(3308) := X"00000000";
		ram_buffer(3309) := X"AF938024";
		ram_buffer(3310) := X"1000FFC4";
		ram_buffer(3311) := X"00000000";
		ram_buffer(3312) := X"27BDFFE0";
		ram_buffer(3313) := X"AFB10018";
		ram_buffer(3314) := X"AFB00014";
		ram_buffer(3315) := X"AFBF001C";
		ram_buffer(3316) := X"00808825";
		ram_buffer(3317) := X"14800005";
		ram_buffer(3318) := X"00A08025";
		ram_buffer(3319) := X"3C040000";
		ram_buffer(3320) := X"24050479";
		ram_buffer(3321) := X"0C00023D";
		ram_buffer(3322) := X"248445CC";
		ram_buffer(3323) := X"16000004";
		ram_buffer(3324) := X"2405047A";
		ram_buffer(3325) := X"3C040000";
		ram_buffer(3326) := X"0C00023D";
		ram_buffer(3327) := X"248445CC";
		ram_buffer(3328) := X"8F828010";
		ram_buffer(3329) := X"00000000";
		ram_buffer(3330) := X"10400004";
		ram_buffer(3331) := X"3C040000";
		ram_buffer(3332) := X"2405047B";
		ram_buffer(3333) := X"0C00023D";
		ram_buffer(3334) := X"248445CC";
		ram_buffer(3335) := X"0C0007DC";
		ram_buffer(3336) := X"00000000";
		ram_buffer(3337) := X"8E230000";
		ram_buffer(3338) := X"8F848034";
		ram_buffer(3339) := X"02038021";
		ram_buffer(3340) := X"0083282B";
		ram_buffer(3341) := X"10A00005";
		ram_buffer(3342) := X"0203182B";
		ram_buffer(3343) := X"10600005";
		ram_buffer(3344) := X"00002825";
		ram_buffer(3345) := X"10000003";
		ram_buffer(3346) := X"0090282B";
		ram_buffer(3347) := X"1060FFFD";
		ram_buffer(3348) := X"24050001";
		ram_buffer(3349) := X"10A00004";
		ram_buffer(3350) := X"AE300000";
		ram_buffer(3351) := X"00002825";
		ram_buffer(3352) := X"0C00075E";
		ram_buffer(3353) := X"02042023";
		ram_buffer(3354) := X"0C000C85";
		ram_buffer(3355) := X"00000000";
		ram_buffer(3356) := X"14400006";
		ram_buffer(3357) := X"00000000";
		ram_buffer(3358) := X"8FBF001C";
		ram_buffer(3359) := X"8FB10018";
		ram_buffer(3360) := X"8FB00014";
		ram_buffer(3361) := X"0800017D";
		ram_buffer(3362) := X"27BD0020";
		ram_buffer(3363) := X"8FBF001C";
		ram_buffer(3364) := X"8FB10018";
		ram_buffer(3365) := X"8FB00014";
		ram_buffer(3366) := X"03E00008";
		ram_buffer(3367) := X"27BD0020";
		ram_buffer(3368) := X"14800007";
		ram_buffer(3369) := X"00000000";
		ram_buffer(3370) := X"0800017D";
		ram_buffer(3371) := X"00000000";
		ram_buffer(3372) := X"8FBF0014";
		ram_buffer(3373) := X"8FB00010";
		ram_buffer(3374) := X"1000FFFB";
		ram_buffer(3375) := X"27BD0018";
		ram_buffer(3376) := X"8F828010";
		ram_buffer(3377) := X"27BDFFE8";
		ram_buffer(3378) := X"AFB00010";
		ram_buffer(3379) := X"AFBF0014";
		ram_buffer(3380) := X"10400005";
		ram_buffer(3381) := X"00808025";
		ram_buffer(3382) := X"3C040000";
		ram_buffer(3383) := X"240504D6";
		ram_buffer(3384) := X"0C00023D";
		ram_buffer(3385) := X"248445CC";
		ram_buffer(3386) := X"0C0007DC";
		ram_buffer(3387) := X"00002825";
		ram_buffer(3388) := X"0C00075E";
		ram_buffer(3389) := X"02002025";
		ram_buffer(3390) := X"0C000C85";
		ram_buffer(3391) := X"00000000";
		ram_buffer(3392) := X"1040FFEB";
		ram_buffer(3393) := X"00000000";
		ram_buffer(3394) := X"8FBF0014";
		ram_buffer(3395) := X"8FB00010";
		ram_buffer(3396) := X"03E00008";
		ram_buffer(3397) := X"27BD0018";
		ram_buffer(3398) := X"27BDFFE0";
		ram_buffer(3399) := X"AFB10018";
		ram_buffer(3400) := X"AFBF001C";
		ram_buffer(3401) := X"AFB00014";
		ram_buffer(3402) := X"0C001160";
		ram_buffer(3403) := X"00808825";
		ram_buffer(3404) := X"2C420010";
		ram_buffer(3405) := X"14400004";
		ram_buffer(3406) := X"240508DD";
		ram_buffer(3407) := X"3C040000";
		ram_buffer(3408) := X"0C00023D";
		ram_buffer(3409) := X"248445CC";
		ram_buffer(3410) := X"0C0007DC";
		ram_buffer(3411) := X"3C0D0000";
		ram_buffer(3412) := X"00006025";
		ram_buffer(3413) := X"25AD46E4";
		ram_buffer(3414) := X"240EFF9C";
		ram_buffer(3415) := X"25840050";
		ram_buffer(3416) := X"02202825";
		ram_buffer(3417) := X"0C000706";
		ram_buffer(3418) := X"01A42021";
		ram_buffer(3419) := X"14400019";
		ram_buffer(3420) := X"00408025";
		ram_buffer(3421) := X"258CFFEC";
		ram_buffer(3422) := X"158EFFF9";
		ram_buffer(3423) := X"25840050";
		ram_buffer(3424) := X"8F848044";
		ram_buffer(3425) := X"0C000706";
		ram_buffer(3426) := X"02202825";
		ram_buffer(3427) := X"14400011";
		ram_buffer(3428) := X"00408025";
		ram_buffer(3429) := X"8F848040";
		ram_buffer(3430) := X"0C000706";
		ram_buffer(3431) := X"02202825";
		ram_buffer(3432) := X"1440000C";
		ram_buffer(3433) := X"00408025";
		ram_buffer(3434) := X"3C040000";
		ram_buffer(3435) := X"02202825";
		ram_buffer(3436) := X"0C000706";
		ram_buffer(3437) := X"24844680";
		ram_buffer(3438) := X"14400006";
		ram_buffer(3439) := X"00408025";
		ram_buffer(3440) := X"3C040000";
		ram_buffer(3441) := X"02202825";
		ram_buffer(3442) := X"0C000706";
		ram_buffer(3443) := X"24844694";
		ram_buffer(3444) := X"00408025";
		ram_buffer(3445) := X"0C000C85";
		ram_buffer(3446) := X"00000000";
		ram_buffer(3447) := X"8FBF001C";
		ram_buffer(3448) := X"02001025";
		ram_buffer(3449) := X"8FB10018";
		ram_buffer(3450) := X"8FB00014";
		ram_buffer(3451) := X"03E00008";
		ram_buffer(3452) := X"27BD0020";
		ram_buffer(3453) := X"27BDFFD8";
		ram_buffer(3454) := X"AFB10018";
		ram_buffer(3455) := X"3C110000";
		ram_buffer(3456) := X"AFB30020";
		ram_buffer(3457) := X"AFB2001C";
		ram_buffer(3458) := X"AFBF0024";
		ram_buffer(3459) := X"AFB00014";
		ram_buffer(3460) := X"26334694";
		ram_buffer(3461) := X"3C120000";
		ram_buffer(3462) := X"8F82803C";
		ram_buffer(3463) := X"00000000";
		ram_buffer(3464) := X"1440000A";
		ram_buffer(3465) := X"00000000";
		ram_buffer(3466) := X"8E4246E4";
		ram_buffer(3467) := X"00000000";
		ram_buffer(3468) := X"2C420002";
		ram_buffer(3469) := X"1440FFF8";
		ram_buffer(3470) := X"00000000";
		ram_buffer(3471) := X"0C00017D";
		ram_buffer(3472) := X"00000000";
		ram_buffer(3473) := X"1000FFF4";
		ram_buffer(3474) := X"00000000";
		ram_buffer(3475) := X"0C0007DC";
		ram_buffer(3476) := X"00000000";
		ram_buffer(3477) := X"8E304694";
		ram_buffer(3478) := X"0C000C85";
		ram_buffer(3479) := X"00000000";
		ram_buffer(3480) := X"1200FFED";
		ram_buffer(3481) := X"00000000";
		ram_buffer(3482) := X"0C000A17";
		ram_buffer(3483) := X"00000000";
		ram_buffer(3484) := X"8E62000C";
		ram_buffer(3485) := X"00000000";
		ram_buffer(3486) := X"8C50000C";
		ram_buffer(3487) := X"0C000289";
		ram_buffer(3488) := X"26040004";
		ram_buffer(3489) := X"8F828038";
		ram_buffer(3490) := X"00000000";
		ram_buffer(3491) := X"2442FFFF";
		ram_buffer(3492) := X"AF828038";
		ram_buffer(3493) := X"8F82803C";
		ram_buffer(3494) := X"00000000";
		ram_buffer(3495) := X"2442FFFF";
		ram_buffer(3496) := X"AF82803C";
		ram_buffer(3497) := X"0C000A2A";
		ram_buffer(3498) := X"00000000";
		ram_buffer(3499) := X"8E040030";
		ram_buffer(3500) := X"0C001030";
		ram_buffer(3501) := X"00000000";
		ram_buffer(3502) := X"0C001030";
		ram_buffer(3503) := X"02002025";
		ram_buffer(3504) := X"1000FFD5";
		ram_buffer(3505) := X"00000000";
		ram_buffer(3506) := X"27BDFFE0";
		ram_buffer(3507) := X"AFB00014";
		ram_buffer(3508) := X"AFBF001C";
		ram_buffer(3509) := X"AFB10018";
		ram_buffer(3510) := X"14800005";
		ram_buffer(3511) := X"00808025";
		ram_buffer(3512) := X"3C040000";
		ram_buffer(3513) := X"24050987";
		ram_buffer(3514) := X"0C00023D";
		ram_buffer(3515) := X"248445CC";
		ram_buffer(3516) := X"0C0007DC";
		ram_buffer(3517) := X"02002025";
		ram_buffer(3518) := X"0C000B70";
		ram_buffer(3519) := X"00000000";
		ram_buffer(3520) := X"24030002";
		ram_buffer(3521) := X"14430026";
		ram_buffer(3522) := X"26110004";
		ram_buffer(3523) := X"0C000289";
		ram_buffer(3524) := X"02202025";
		ram_buffer(3525) := X"0C000A17";
		ram_buffer(3526) := X"00000000";
		ram_buffer(3527) := X"8E020028";
		ram_buffer(3528) := X"00000000";
		ram_buffer(3529) := X"10400005";
		ram_buffer(3530) := X"00000000";
		ram_buffer(3531) := X"0C000289";
		ram_buffer(3532) := X"26040018";
		ram_buffer(3533) := X"24020001";
		ram_buffer(3534) := X"A2020055";
		ram_buffer(3535) := X"0C000A2A";
		ram_buffer(3536) := X"00000000";
		ram_buffer(3537) := X"8E04002C";
		ram_buffer(3538) := X"8F828030";
		ram_buffer(3539) := X"00000000";
		ram_buffer(3540) := X"0044102B";
		ram_buffer(3541) := X"10400003";
		ram_buffer(3542) := X"00041080";
		ram_buffer(3543) := X"AF848030";
		ram_buffer(3544) := X"00041080";
		ram_buffer(3545) := X"00441021";
		ram_buffer(3546) := X"3C040000";
		ram_buffer(3547) := X"00021080";
		ram_buffer(3548) := X"248446E4";
		ram_buffer(3549) := X"00822021";
		ram_buffer(3550) := X"0C000260";
		ram_buffer(3551) := X"02202825";
		ram_buffer(3552) := X"8F83800C";
		ram_buffer(3553) := X"8E02002C";
		ram_buffer(3554) := X"8C63002C";
		ram_buffer(3555) := X"00000000";
		ram_buffer(3556) := X"0062102B";
		ram_buffer(3557) := X"10400002";
		ram_buffer(3558) := X"24020001";
		ram_buffer(3559) := X"AF828024";
		ram_buffer(3560) := X"0C000C85";
		ram_buffer(3561) := X"00000000";
		ram_buffer(3562) := X"8FBF001C";
		ram_buffer(3563) := X"8FB10018";
		ram_buffer(3564) := X"8FB00014";
		ram_buffer(3565) := X"00001025";
		ram_buffer(3566) := X"03E00008";
		ram_buffer(3567) := X"27BD0020";
		ram_buffer(3568) := X"27BDFFE0";
		ram_buffer(3569) := X"AFB20018";
		ram_buffer(3570) := X"AFB10014";
		ram_buffer(3571) := X"AFBF001C";
		ram_buffer(3572) := X"AFB00010";
		ram_buffer(3573) := X"00808825";
		ram_buffer(3574) := X"14800005";
		ram_buffer(3575) := X"00A09025";
		ram_buffer(3576) := X"3C040000";
		ram_buffer(3577) := X"24050BDA";
		ram_buffer(3578) := X"0C00023D";
		ram_buffer(3579) := X"248445CC";
		ram_buffer(3580) := X"16400004";
		ram_buffer(3581) := X"3C040000";
		ram_buffer(3582) := X"24050BDB";
		ram_buffer(3583) := X"0C00023D";
		ram_buffer(3584) := X"248445CC";
		ram_buffer(3585) := X"0C000A17";
		ram_buffer(3586) := X"00000000";
		ram_buffer(3587) := X"8F848034";
		ram_buffer(3588) := X"8F82800C";
		ram_buffer(3589) := X"00000000";
		ram_buffer(3590) := X"90420055";
		ram_buffer(3591) := X"00000000";
		ram_buffer(3592) := X"1040000D";
		ram_buffer(3593) := X"2402FFFF";
		ram_buffer(3594) := X"8F82800C";
		ram_buffer(3595) := X"24100001";
		ram_buffer(3596) := X"A0400055";
		ram_buffer(3597) := X"0C000A2A";
		ram_buffer(3598) := X"00000000";
		ram_buffer(3599) := X"8FBF001C";
		ram_buffer(3600) := X"02001025";
		ram_buffer(3601) := X"8FB20018";
		ram_buffer(3602) := X"8FB10014";
		ram_buffer(3603) := X"8FB00010";
		ram_buffer(3604) := X"03E00008";
		ram_buffer(3605) := X"27BD0020";
		ram_buffer(3606) := X"8E430000";
		ram_buffer(3607) := X"00000000";
		ram_buffer(3608) := X"1062FFF4";
		ram_buffer(3609) := X"00008025";
		ram_buffer(3610) := X"8F858020";
		ram_buffer(3611) := X"8E260000";
		ram_buffer(3612) := X"8E220004";
		ram_buffer(3613) := X"10C50003";
		ram_buffer(3614) := X"0082282B";
		ram_buffer(3615) := X"10A0FFED";
		ram_buffer(3616) := X"24100001";
		ram_buffer(3617) := X"00822823";
		ram_buffer(3618) := X"00A3282B";
		ram_buffer(3619) := X"10A0FFE9";
		ram_buffer(3620) := X"24100001";
		ram_buffer(3621) := X"00641823";
		ram_buffer(3622) := X"00621821";
		ram_buffer(3623) := X"AE430000";
		ram_buffer(3624) := X"0C000968";
		ram_buffer(3625) := X"02202025";
		ram_buffer(3626) := X"1000FFE2";
		ram_buffer(3627) := X"00008025";
		ram_buffer(3628) := X"8F82800C";
		ram_buffer(3629) := X"8F84800C";
		ram_buffer(3630) := X"8F83800C";
		ram_buffer(3631) := X"8C420018";
		ram_buffer(3632) := X"8C65002C";
		ram_buffer(3633) := X"24030005";
		ram_buffer(3634) := X"00651823";
		ram_buffer(3635) := X"03E00008";
		ram_buffer(3636) := X"AC830018";
		ram_buffer(3637) := X"8F82800C";
		ram_buffer(3638) := X"00000000";
		ram_buffer(3639) := X"10400007";
		ram_buffer(3640) := X"00000000";
		ram_buffer(3641) := X"8F83800C";
		ram_buffer(3642) := X"00000000";
		ram_buffer(3643) := X"8C62004C";
		ram_buffer(3644) := X"00000000";
		ram_buffer(3645) := X"24420001";
		ram_buffer(3646) := X"AC62004C";
		ram_buffer(3647) := X"8F82800C";
		ram_buffer(3648) := X"03E00008";
		ram_buffer(3649) := X"00000000";
		ram_buffer(3650) := X"27BDFFE0";
		ram_buffer(3651) := X"AFB10018";
		ram_buffer(3652) := X"AFB00014";
		ram_buffer(3653) := X"AFBF001C";
		ram_buffer(3654) := X"00808825";
		ram_buffer(3655) := X"0C000A17";
		ram_buffer(3656) := X"00A08025";
		ram_buffer(3657) := X"8F82800C";
		ram_buffer(3658) := X"00000000";
		ram_buffer(3659) := X"8C420050";
		ram_buffer(3660) := X"00000000";
		ram_buffer(3661) := X"1440000A";
		ram_buffer(3662) := X"00000000";
		ram_buffer(3663) := X"8F82800C";
		ram_buffer(3664) := X"24030001";
		ram_buffer(3665) := X"A0430054";
		ram_buffer(3666) := X"12000005";
		ram_buffer(3667) := X"24050001";
		ram_buffer(3668) := X"0C00075E";
		ram_buffer(3669) := X"02002025";
		ram_buffer(3670) := X"0C00017D";
		ram_buffer(3671) := X"00000000";
		ram_buffer(3672) := X"0C000A2A";
		ram_buffer(3673) := X"00000000";
		ram_buffer(3674) := X"0C000A17";
		ram_buffer(3675) := X"00000000";
		ram_buffer(3676) := X"8F82800C";
		ram_buffer(3677) := X"00000000";
		ram_buffer(3678) := X"8C500050";
		ram_buffer(3679) := X"00000000";
		ram_buffer(3680) := X"12000005";
		ram_buffer(3681) := X"00000000";
		ram_buffer(3682) := X"8F82800C";
		ram_buffer(3683) := X"1220000D";
		ram_buffer(3684) := X"2603FFFF";
		ram_buffer(3685) := X"AC400050";
		ram_buffer(3686) := X"8F82800C";
		ram_buffer(3687) := X"00000000";
		ram_buffer(3688) := X"A0400054";
		ram_buffer(3689) := X"0C000A2A";
		ram_buffer(3690) := X"00000000";
		ram_buffer(3691) := X"8FBF001C";
		ram_buffer(3692) := X"02001025";
		ram_buffer(3693) := X"8FB10018";
		ram_buffer(3694) := X"8FB00014";
		ram_buffer(3695) := X"03E00008";
		ram_buffer(3696) := X"27BD0020";
		ram_buffer(3697) := X"AC430050";
		ram_buffer(3698) := X"1000FFF3";
		ram_buffer(3699) := X"00000000";
		ram_buffer(3700) := X"27BDFFD8";
		ram_buffer(3701) := X"AFB30020";
		ram_buffer(3702) := X"AFB2001C";
		ram_buffer(3703) := X"AFB10018";
		ram_buffer(3704) := X"AFB00014";
		ram_buffer(3705) := X"AFBF0024";
		ram_buffer(3706) := X"00808825";
		ram_buffer(3707) := X"00A08025";
		ram_buffer(3708) := X"00C09025";
		ram_buffer(3709) := X"0C000A17";
		ram_buffer(3710) := X"00E09825";
		ram_buffer(3711) := X"8F82800C";
		ram_buffer(3712) := X"24030002";
		ram_buffer(3713) := X"90420054";
		ram_buffer(3714) := X"00000000";
		ram_buffer(3715) := X"304200FF";
		ram_buffer(3716) := X"10430010";
		ram_buffer(3717) := X"00000000";
		ram_buffer(3718) := X"8F82800C";
		ram_buffer(3719) := X"00118827";
		ram_buffer(3720) := X"8C440050";
		ram_buffer(3721) := X"24030001";
		ram_buffer(3722) := X"02248824";
		ram_buffer(3723) := X"AC510050";
		ram_buffer(3724) := X"8F82800C";
		ram_buffer(3725) := X"00000000";
		ram_buffer(3726) := X"A0430054";
		ram_buffer(3727) := X"12600005";
		ram_buffer(3728) := X"24050001";
		ram_buffer(3729) := X"0C00075E";
		ram_buffer(3730) := X"02602025";
		ram_buffer(3731) := X"0C00017D";
		ram_buffer(3732) := X"00000000";
		ram_buffer(3733) := X"0C000A2A";
		ram_buffer(3734) := X"00000000";
		ram_buffer(3735) := X"0C000A17";
		ram_buffer(3736) := X"00000000";
		ram_buffer(3737) := X"12400006";
		ram_buffer(3738) := X"00000000";
		ram_buffer(3739) := X"8F82800C";
		ram_buffer(3740) := X"00000000";
		ram_buffer(3741) := X"8C420050";
		ram_buffer(3742) := X"00000000";
		ram_buffer(3743) := X"AE420000";
		ram_buffer(3744) := X"8F82800C";
		ram_buffer(3745) := X"00008825";
		ram_buffer(3746) := X"90430054";
		ram_buffer(3747) := X"24020001";
		ram_buffer(3748) := X"306300FF";
		ram_buffer(3749) := X"10620007";
		ram_buffer(3750) := X"00000000";
		ram_buffer(3751) := X"8F82800C";
		ram_buffer(3752) := X"00108027";
		ram_buffer(3753) := X"8C430050";
		ram_buffer(3754) := X"24110001";
		ram_buffer(3755) := X"02038024";
		ram_buffer(3756) := X"AC500050";
		ram_buffer(3757) := X"8F82800C";
		ram_buffer(3758) := X"00000000";
		ram_buffer(3759) := X"A0400054";
		ram_buffer(3760) := X"0C000A2A";
		ram_buffer(3761) := X"00000000";
		ram_buffer(3762) := X"8FBF0024";
		ram_buffer(3763) := X"02201025";
		ram_buffer(3764) := X"8FB30020";
		ram_buffer(3765) := X"8FB2001C";
		ram_buffer(3766) := X"8FB10018";
		ram_buffer(3767) := X"8FB00014";
		ram_buffer(3768) := X"03E00008";
		ram_buffer(3769) := X"27BD0028";
		ram_buffer(3770) := X"27BDFFD8";
		ram_buffer(3771) := X"AFB30020";
		ram_buffer(3772) := X"AFB2001C";
		ram_buffer(3773) := X"AFB10018";
		ram_buffer(3774) := X"AFB00014";
		ram_buffer(3775) := X"AFBF0024";
		ram_buffer(3776) := X"00808025";
		ram_buffer(3777) := X"00A09025";
		ram_buffer(3778) := X"00C08825";
		ram_buffer(3779) := X"14800005";
		ram_buffer(3780) := X"00E09825";
		ram_buffer(3781) := X"3C040000";
		ram_buffer(3782) := X"2405110C";
		ram_buffer(3783) := X"0C00023D";
		ram_buffer(3784) := X"248445CC";
		ram_buffer(3785) := X"0C000A17";
		ram_buffer(3786) := X"00000000";
		ram_buffer(3787) := X"12600004";
		ram_buffer(3788) := X"00000000";
		ram_buffer(3789) := X"8E020050";
		ram_buffer(3790) := X"00000000";
		ram_buffer(3791) := X"AE620000";
		ram_buffer(3792) := X"92030054";
		ram_buffer(3793) := X"24020002";
		ram_buffer(3794) := X"A2020054";
		ram_buffer(3795) := X"24020002";
		ram_buffer(3796) := X"12220023";
		ram_buffer(3797) := X"306300FF";
		ram_buffer(3798) := X"2E240003";
		ram_buffer(3799) := X"10800009";
		ram_buffer(3800) := X"00000000";
		ram_buffer(3801) := X"24020001";
		ram_buffer(3802) := X"12220017";
		ram_buffer(3803) := X"00000000";
		ram_buffer(3804) := X"24020001";
		ram_buffer(3805) := X"10620020";
		ram_buffer(3806) := X"00000000";
		ram_buffer(3807) := X"10000008";
		ram_buffer(3808) := X"24110001";
		ram_buffer(3809) := X"24040003";
		ram_buffer(3810) := X"12240012";
		ram_buffer(3811) := X"24040004";
		ram_buffer(3812) := X"1624FFF7";
		ram_buffer(3813) := X"00000000";
		ram_buffer(3814) := X"1462000E";
		ram_buffer(3815) := X"00008825";
		ram_buffer(3816) := X"0C000A2A";
		ram_buffer(3817) := X"00000000";
		ram_buffer(3818) := X"8FBF0024";
		ram_buffer(3819) := X"02201025";
		ram_buffer(3820) := X"8FB30020";
		ram_buffer(3821) := X"8FB2001C";
		ram_buffer(3822) := X"8FB10018";
		ram_buffer(3823) := X"8FB00014";
		ram_buffer(3824) := X"03E00008";
		ram_buffer(3825) := X"27BD0028";
		ram_buffer(3826) := X"8E020050";
		ram_buffer(3827) := X"00000000";
		ram_buffer(3828) := X"00529025";
		ram_buffer(3829) := X"AE120050";
		ram_buffer(3830) := X"1000FFE6";
		ram_buffer(3831) := X"24020001";
		ram_buffer(3832) := X"8E020050";
		ram_buffer(3833) := X"00000000";
		ram_buffer(3834) := X"24420001";
		ram_buffer(3835) := X"AE020050";
		ram_buffer(3836) := X"1000FFE0";
		ram_buffer(3837) := X"24020001";
		ram_buffer(3838) := X"26110004";
		ram_buffer(3839) := X"0C000289";
		ram_buffer(3840) := X"02202025";
		ram_buffer(3841) := X"8E04002C";
		ram_buffer(3842) := X"8F828030";
		ram_buffer(3843) := X"00000000";
		ram_buffer(3844) := X"0044102B";
		ram_buffer(3845) := X"10400003";
		ram_buffer(3846) := X"00041080";
		ram_buffer(3847) := X"AF848030";
		ram_buffer(3848) := X"00041080";
		ram_buffer(3849) := X"00441021";
		ram_buffer(3850) := X"3C040000";
		ram_buffer(3851) := X"00021080";
		ram_buffer(3852) := X"248446E4";
		ram_buffer(3853) := X"00822021";
		ram_buffer(3854) := X"0C000260";
		ram_buffer(3855) := X"02202825";
		ram_buffer(3856) := X"8E020028";
		ram_buffer(3857) := X"00000000";
		ram_buffer(3858) := X"10400004";
		ram_buffer(3859) := X"3C040000";
		ram_buffer(3860) := X"24051144";
		ram_buffer(3861) := X"0C00023D";
		ram_buffer(3862) := X"248445CC";
		ram_buffer(3863) := X"8F83800C";
		ram_buffer(3864) := X"8E02002C";
		ram_buffer(3865) := X"8C63002C";
		ram_buffer(3866) := X"00000000";
		ram_buffer(3867) := X"0062102B";
		ram_buffer(3868) := X"1040FFC2";
		ram_buffer(3869) := X"00000000";
		ram_buffer(3870) := X"0C00017D";
		ram_buffer(3871) := X"24110001";
		ram_buffer(3872) := X"1000FFC7";
		ram_buffer(3873) := X"00000000";
		ram_buffer(3874) := X"27BDFFD8";
		ram_buffer(3875) := X"AFB40020";
		ram_buffer(3876) := X"AFB3001C";
		ram_buffer(3877) := X"AFB20018";
		ram_buffer(3878) := X"AFB10014";
		ram_buffer(3879) := X"AFB00010";
		ram_buffer(3880) := X"AFBF0024";
		ram_buffer(3881) := X"00808025";
		ram_buffer(3882) := X"00A09825";
		ram_buffer(3883) := X"00C08825";
		ram_buffer(3884) := X"8FB20038";
		ram_buffer(3885) := X"14800005";
		ram_buffer(3886) := X"00E0A025";
		ram_buffer(3887) := X"3C040000";
		ram_buffer(3888) := X"24051177";
		ram_buffer(3889) := X"0C00023D";
		ram_buffer(3890) := X"248445CC";
		ram_buffer(3891) := X"12800004";
		ram_buffer(3892) := X"00000000";
		ram_buffer(3893) := X"8E020050";
		ram_buffer(3894) := X"00000000";
		ram_buffer(3895) := X"AE820000";
		ram_buffer(3896) := X"92030054";
		ram_buffer(3897) := X"24020002";
		ram_buffer(3898) := X"24040002";
		ram_buffer(3899) := X"306300FF";
		ram_buffer(3900) := X"A2020054";
		ram_buffer(3901) := X"12240021";
		ram_buffer(3902) := X"00000000";
		ram_buffer(3903) := X"2E220003";
		ram_buffer(3904) := X"10400009";
		ram_buffer(3905) := X"24020003";
		ram_buffer(3906) := X"24020001";
		ram_buffer(3907) := X"12220015";
		ram_buffer(3908) := X"00000000";
		ram_buffer(3909) := X"24020001";
		ram_buffer(3910) := X"1062001E";
		ram_buffer(3911) := X"00000000";
		ram_buffer(3912) := X"10000008";
		ram_buffer(3913) := X"24020001";
		ram_buffer(3914) := X"12220011";
		ram_buffer(3915) := X"00000000";
		ram_buffer(3916) := X"24020004";
		ram_buffer(3917) := X"1622FFF7";
		ram_buffer(3918) := X"00000000";
		ram_buffer(3919) := X"1464000C";
		ram_buffer(3920) := X"00001025";
		ram_buffer(3921) := X"8FBF0024";
		ram_buffer(3922) := X"8FB40020";
		ram_buffer(3923) := X"8FB3001C";
		ram_buffer(3924) := X"8FB20018";
		ram_buffer(3925) := X"8FB10014";
		ram_buffer(3926) := X"8FB00010";
		ram_buffer(3927) := X"03E00008";
		ram_buffer(3928) := X"27BD0028";
		ram_buffer(3929) := X"8E020050";
		ram_buffer(3930) := X"00000000";
		ram_buffer(3931) := X"00539825";
		ram_buffer(3932) := X"AE130050";
		ram_buffer(3933) := X"1000FFE8";
		ram_buffer(3934) := X"24020001";
		ram_buffer(3935) := X"8E020050";
		ram_buffer(3936) := X"00000000";
		ram_buffer(3937) := X"24420001";
		ram_buffer(3938) := X"AE020050";
		ram_buffer(3939) := X"1000FFE2";
		ram_buffer(3940) := X"24020001";
		ram_buffer(3941) := X"8E020028";
		ram_buffer(3942) := X"00000000";
		ram_buffer(3943) := X"10400004";
		ram_buffer(3944) := X"240511BE";
		ram_buffer(3945) := X"3C040000";
		ram_buffer(3946) := X"0C00023D";
		ram_buffer(3947) := X"248445CC";
		ram_buffer(3948) := X"8F828010";
		ram_buffer(3949) := X"00000000";
		ram_buffer(3950) := X"1440001F";
		ram_buffer(3951) := X"3C040000";
		ram_buffer(3952) := X"26110004";
		ram_buffer(3953) := X"0C000289";
		ram_buffer(3954) := X"02202025";
		ram_buffer(3955) := X"8E04002C";
		ram_buffer(3956) := X"8F828030";
		ram_buffer(3957) := X"00000000";
		ram_buffer(3958) := X"0044102B";
		ram_buffer(3959) := X"10400003";
		ram_buffer(3960) := X"00041080";
		ram_buffer(3961) := X"AF848030";
		ram_buffer(3962) := X"00041080";
		ram_buffer(3963) := X"00441021";
		ram_buffer(3964) := X"3C040000";
		ram_buffer(3965) := X"00021080";
		ram_buffer(3966) := X"248446E4";
		ram_buffer(3967) := X"02202825";
		ram_buffer(3968) := X"00822021";
		ram_buffer(3969) := X"0C000260";
		ram_buffer(3970) := X"00000000";
		ram_buffer(3971) := X"8F83800C";
		ram_buffer(3972) := X"8E02002C";
		ram_buffer(3973) := X"8C63002C";
		ram_buffer(3974) := X"00000000";
		ram_buffer(3975) := X"0062102B";
		ram_buffer(3976) := X"1040FFBF";
		ram_buffer(3977) := X"00000000";
		ram_buffer(3978) := X"12400006";
		ram_buffer(3979) := X"24020001";
		ram_buffer(3980) := X"1000FFC4";
		ram_buffer(3981) := X"AE420000";
		ram_buffer(3982) := X"26050018";
		ram_buffer(3983) := X"1000FFF1";
		ram_buffer(3984) := X"248446A8";
		ram_buffer(3985) := X"AF828024";
		ram_buffer(3986) := X"1000FFBE";
		ram_buffer(3987) := X"00000000";
		ram_buffer(3988) := X"27BDFFE0";
		ram_buffer(3989) := X"AFB10014";
		ram_buffer(3990) := X"AFB00010";
		ram_buffer(3991) := X"AFBF001C";
		ram_buffer(3992) := X"AFB20018";
		ram_buffer(3993) := X"00808025";
		ram_buffer(3994) := X"14800005";
		ram_buffer(3995) := X"00A08825";
		ram_buffer(3996) := X"3C040000";
		ram_buffer(3997) := X"240511F2";
		ram_buffer(3998) := X"0C00023D";
		ram_buffer(3999) := X"248445CC";
		ram_buffer(4000) := X"24030002";
		ram_buffer(4001) := X"92020054";
		ram_buffer(4002) := X"A2030054";
		ram_buffer(4003) := X"8E030050";
		ram_buffer(4004) := X"304200FF";
		ram_buffer(4005) := X"24630001";
		ram_buffer(4006) := X"AE030050";
		ram_buffer(4007) := X"24030001";
		ram_buffer(4008) := X"14430029";
		ram_buffer(4009) := X"00000000";
		ram_buffer(4010) := X"8E020028";
		ram_buffer(4011) := X"00000000";
		ram_buffer(4012) := X"10400004";
		ram_buffer(4013) := X"24051218";
		ram_buffer(4014) := X"3C040000";
		ram_buffer(4015) := X"0C00023D";
		ram_buffer(4016) := X"248445CC";
		ram_buffer(4017) := X"8F828010";
		ram_buffer(4018) := X"00000000";
		ram_buffer(4019) := X"14400024";
		ram_buffer(4020) := X"3C040000";
		ram_buffer(4021) := X"26120004";
		ram_buffer(4022) := X"0C000289";
		ram_buffer(4023) := X"02402025";
		ram_buffer(4024) := X"8E04002C";
		ram_buffer(4025) := X"8F828030";
		ram_buffer(4026) := X"00000000";
		ram_buffer(4027) := X"0044102B";
		ram_buffer(4028) := X"10400003";
		ram_buffer(4029) := X"00041080";
		ram_buffer(4030) := X"AF848030";
		ram_buffer(4031) := X"00041080";
		ram_buffer(4032) := X"00441021";
		ram_buffer(4033) := X"3C040000";
		ram_buffer(4034) := X"00021080";
		ram_buffer(4035) := X"248446E4";
		ram_buffer(4036) := X"02402825";
		ram_buffer(4037) := X"00822021";
		ram_buffer(4038) := X"0C000260";
		ram_buffer(4039) := X"00000000";
		ram_buffer(4040) := X"8F83800C";
		ram_buffer(4041) := X"8E02002C";
		ram_buffer(4042) := X"8C63002C";
		ram_buffer(4043) := X"00000000";
		ram_buffer(4044) := X"0062102B";
		ram_buffer(4045) := X"10400004";
		ram_buffer(4046) := X"00000000";
		ram_buffer(4047) := X"1220000B";
		ram_buffer(4048) := X"24020001";
		ram_buffer(4049) := X"AE220000";
		ram_buffer(4050) := X"8FBF001C";
		ram_buffer(4051) := X"8FB20018";
		ram_buffer(4052) := X"8FB10014";
		ram_buffer(4053) := X"8FB00010";
		ram_buffer(4054) := X"03E00008";
		ram_buffer(4055) := X"27BD0020";
		ram_buffer(4056) := X"26050018";
		ram_buffer(4057) := X"1000FFEC";
		ram_buffer(4058) := X"248446A8";
		ram_buffer(4059) := X"AF828024";
		ram_buffer(4060) := X"1000FFF5";
		ram_buffer(4061) := X"00000000";
		ram_buffer(4062) := X"27BDFFE0";
		ram_buffer(4063) := X"AFB00014";
		ram_buffer(4064) := X"AFBF001C";
		ram_buffer(4065) := X"AFB10018";
		ram_buffer(4066) := X"14800002";
		ram_buffer(4067) := X"00808025";
		ram_buffer(4068) := X"8F90800C";
		ram_buffer(4069) := X"0C000A17";
		ram_buffer(4070) := X"00000000";
		ram_buffer(4071) := X"92030054";
		ram_buffer(4072) := X"24020002";
		ram_buffer(4073) := X"306300FF";
		ram_buffer(4074) := X"14620003";
		ram_buffer(4075) := X"00008825";
		ram_buffer(4076) := X"A2000054";
		ram_buffer(4077) := X"24110001";
		ram_buffer(4078) := X"0C000A2A";
		ram_buffer(4079) := X"00000000";
		ram_buffer(4080) := X"8FBF001C";
		ram_buffer(4081) := X"02201025";
		ram_buffer(4082) := X"8FB00014";
		ram_buffer(4083) := X"8FB10018";
		ram_buffer(4084) := X"03E00008";
		ram_buffer(4085) := X"27BD0020";
		ram_buffer(4086) := X"03E00008";
		ram_buffer(4087) := X"00000000";
		ram_buffer(4088) := X"27BDFFE8";
		ram_buffer(4089) := X"AFBF0014";
		ram_buffer(4090) := X"0C00014C";
		ram_buffer(4091) := X"00000000";
		ram_buffer(4092) := X"0C000233";
		ram_buffer(4093) := X"00000000";
		ram_buffer(4094) := X"0C00015B";
		ram_buffer(4095) := X"00000000";
		ram_buffer(4096) := X"0C000238";
		ram_buffer(4097) := X"00000000";
		ram_buffer(4098) := X"1000FFFF";
		ram_buffer(4099) := X"00000000";
		ram_buffer(4100) := X"3C040000";
		ram_buffer(4101) := X"24050070";
		ram_buffer(4102) := X"0800023D";
		ram_buffer(4103) := X"248445EC";
		ram_buffer(4104) := X"27BDFFE0";
		ram_buffer(4105) := X"30820003";
		ram_buffer(4106) := X"AFB00014";
		ram_buffer(4107) := X"AFBF001C";
		ram_buffer(4108) := X"AFB10018";
		ram_buffer(4109) := X"10400004";
		ram_buffer(4110) := X"00808025";
		ram_buffer(4111) := X"2404FFFC";
		ram_buffer(4112) := X"02048024";
		ram_buffer(4113) := X"26100004";
		ram_buffer(4114) := X"0C0007DC";
		ram_buffer(4115) := X"00000000";
		ram_buffer(4116) := X"8F82804C";
		ram_buffer(4117) := X"00000000";
		ram_buffer(4118) := X"14400005";
		ram_buffer(4119) := X"3C020000";
		ram_buffer(4120) := X"2403FFFC";
		ram_buffer(4121) := X"2442474C";
		ram_buffer(4122) := X"00431024";
		ram_buffer(4123) := X"AF82804C";
		ram_buffer(4124) := X"8F828050";
		ram_buffer(4125) := X"00000000";
		ram_buffer(4126) := X"02028021";
		ram_buffer(4127) := X"2E031FFC";
		ram_buffer(4128) := X"10600007";
		ram_buffer(4129) := X"00008825";
		ram_buffer(4130) := X"0050182B";
		ram_buffer(4131) := X"10600004";
		ram_buffer(4132) := X"00000000";
		ram_buffer(4133) := X"8F91804C";
		ram_buffer(4134) := X"AF908050";
		ram_buffer(4135) := X"02228821";
		ram_buffer(4136) := X"0C000C85";
		ram_buffer(4137) := X"00000000";
		ram_buffer(4138) := X"8FBF001C";
		ram_buffer(4139) := X"02201025";
		ram_buffer(4140) := X"8FB00014";
		ram_buffer(4141) := X"8FB10018";
		ram_buffer(4142) := X"03E00008";
		ram_buffer(4143) := X"27BD0020";
		ram_buffer(4144) := X"10800004";
		ram_buffer(4145) := X"3C040000";
		ram_buffer(4146) := X"240500AB";
		ram_buffer(4147) := X"0800023D";
		ram_buffer(4148) := X"24844604";
		ram_buffer(4149) := X"03E00008";
		ram_buffer(4150) := X"00000000";
		ram_buffer(4151) := X"03E00008";
		ram_buffer(4152) := X"AF808050";
		ram_buffer(4153) := X"8F828050";
		ram_buffer(4154) := X"24031FFC";
		ram_buffer(4155) := X"03E00008";
		ram_buffer(4156) := X"00621023";
		ram_buffer(4157) := X"28CA0008";
		ram_buffer(4158) := X"1540005B";
		ram_buffer(4159) := X"00801025";
		ram_buffer(4160) := X"00A4C026";
		ram_buffer(4161) := X"33180003";
		ram_buffer(4162) := X"17000066";
		ram_buffer(4163) := X"00043823";
		ram_buffer(4164) := X"30E70003";
		ram_buffer(4165) := X"10E00005";
		ram_buffer(4166) := X"00C73023";
		ram_buffer(4167) := X"88B80000";
		ram_buffer(4168) := X"00A72821";
		ram_buffer(4169) := X"A8980000";
		ram_buffer(4170) := X"00872021";
		ram_buffer(4171) := X"30D8003F";
		ram_buffer(4172) := X"10D80026";
		ram_buffer(4173) := X"00D83823";
		ram_buffer(4174) := X"00873821";
		ram_buffer(4175) := X"8CA80000";
		ram_buffer(4176) := X"8CA90004";
		ram_buffer(4177) := X"8CAA0008";
		ram_buffer(4178) := X"8CAB000C";
		ram_buffer(4179) := X"8CAC0010";
		ram_buffer(4180) := X"8CAD0014";
		ram_buffer(4181) := X"8CAE0018";
		ram_buffer(4182) := X"8CAF001C";
		ram_buffer(4183) := X"AC880000";
		ram_buffer(4184) := X"AC890004";
		ram_buffer(4185) := X"AC8A0008";
		ram_buffer(4186) := X"AC8B000C";
		ram_buffer(4187) := X"AC8C0010";
		ram_buffer(4188) := X"AC8D0014";
		ram_buffer(4189) := X"AC8E0018";
		ram_buffer(4190) := X"AC8F001C";
		ram_buffer(4191) := X"8CA80020";
		ram_buffer(4192) := X"8CA90024";
		ram_buffer(4193) := X"8CAA0028";
		ram_buffer(4194) := X"8CAB002C";
		ram_buffer(4195) := X"8CAC0030";
		ram_buffer(4196) := X"8CAD0034";
		ram_buffer(4197) := X"8CAE0038";
		ram_buffer(4198) := X"8CAF003C";
		ram_buffer(4199) := X"AC880020";
		ram_buffer(4200) := X"AC890024";
		ram_buffer(4201) := X"AC8A0028";
		ram_buffer(4202) := X"AC8B002C";
		ram_buffer(4203) := X"AC8C0030";
		ram_buffer(4204) := X"AC8D0034";
		ram_buffer(4205) := X"AC8E0038";
		ram_buffer(4206) := X"AC8F003C";
		ram_buffer(4207) := X"24840040";
		ram_buffer(4208) := X"1487FFDE";
		ram_buffer(4209) := X"24A50040";
		ram_buffer(4210) := X"03003025";
		ram_buffer(4211) := X"30D8001F";
		ram_buffer(4212) := X"10D80013";
		ram_buffer(4213) := X"00000000";
		ram_buffer(4214) := X"8CA80000";
		ram_buffer(4215) := X"8CA90004";
		ram_buffer(4216) := X"8CAA0008";
		ram_buffer(4217) := X"8CAB000C";
		ram_buffer(4218) := X"8CAC0010";
		ram_buffer(4219) := X"8CAD0014";
		ram_buffer(4220) := X"8CAE0018";
		ram_buffer(4221) := X"8CAF001C";
		ram_buffer(4222) := X"24A50020";
		ram_buffer(4223) := X"AC880000";
		ram_buffer(4224) := X"AC890004";
		ram_buffer(4225) := X"AC8A0008";
		ram_buffer(4226) := X"AC8B000C";
		ram_buffer(4227) := X"AC8C0010";
		ram_buffer(4228) := X"AC8D0014";
		ram_buffer(4229) := X"AC8E0018";
		ram_buffer(4230) := X"AC8F001C";
		ram_buffer(4231) := X"24840020";
		ram_buffer(4232) := X"33060003";
		ram_buffer(4233) := X"10D80007";
		ram_buffer(4234) := X"03063823";
		ram_buffer(4235) := X"00873821";
		ram_buffer(4236) := X"8CAB0000";
		ram_buffer(4237) := X"24840004";
		ram_buffer(4238) := X"24A50004";
		ram_buffer(4239) := X"1487FFFC";
		ram_buffer(4240) := X"AC8BFFFC";
		ram_buffer(4241) := X"18C00006";
		ram_buffer(4242) := X"00863821";
		ram_buffer(4243) := X"80A30000";
		ram_buffer(4244) := X"24840001";
		ram_buffer(4245) := X"24A50001";
		ram_buffer(4246) := X"1487FFFC";
		ram_buffer(4247) := X"A083FFFF";
		ram_buffer(4248) := X"03E00008";
		ram_buffer(4249) := X"00000000";
		ram_buffer(4250) := X"30D80003";
		ram_buffer(4251) := X"1306FFF5";
		ram_buffer(4252) := X"30990003";
		ram_buffer(4253) := X"1720FFF3";
		ram_buffer(4254) := X"30B90003";
		ram_buffer(4255) := X"1720FFF1";
		ram_buffer(4256) := X"00D83823";
		ram_buffer(4257) := X"00873821";
		ram_buffer(4258) := X"8CAB0000";
		ram_buffer(4259) := X"24840004";
		ram_buffer(4260) := X"24A50004";
		ram_buffer(4261) := X"1487FFFC";
		ram_buffer(4262) := X"AC8BFFFC";
		ram_buffer(4263) := X"1000FFE9";
		ram_buffer(4264) := X"03003025";
		ram_buffer(4265) := X"30E70003";
		ram_buffer(4266) := X"10E00006";
		ram_buffer(4267) := X"00C73023";
		ram_buffer(4268) := X"88A30000";
		ram_buffer(4269) := X"98A30003";
		ram_buffer(4270) := X"00A72821";
		ram_buffer(4271) := X"A8830000";
		ram_buffer(4272) := X"00872021";
		ram_buffer(4273) := X"30D8003F";
		ram_buffer(4274) := X"10D80036";
		ram_buffer(4275) := X"00D83823";
		ram_buffer(4276) := X"00873821";
		ram_buffer(4277) := X"88A80000";
		ram_buffer(4278) := X"88A90004";
		ram_buffer(4279) := X"88AA0008";
		ram_buffer(4280) := X"88AB000C";
		ram_buffer(4281) := X"88AC0010";
		ram_buffer(4282) := X"88AD0014";
		ram_buffer(4283) := X"88AE0018";
		ram_buffer(4284) := X"88AF001C";
		ram_buffer(4285) := X"98A80003";
		ram_buffer(4286) := X"98A90007";
		ram_buffer(4287) := X"98AA000B";
		ram_buffer(4288) := X"98AB000F";
		ram_buffer(4289) := X"98AC0013";
		ram_buffer(4290) := X"98AD0017";
		ram_buffer(4291) := X"98AE001B";
		ram_buffer(4292) := X"98AF001F";
		ram_buffer(4293) := X"AC880000";
		ram_buffer(4294) := X"AC890004";
		ram_buffer(4295) := X"AC8A0008";
		ram_buffer(4296) := X"AC8B000C";
		ram_buffer(4297) := X"AC8C0010";
		ram_buffer(4298) := X"AC8D0014";
		ram_buffer(4299) := X"AC8E0018";
		ram_buffer(4300) := X"AC8F001C";
		ram_buffer(4301) := X"88A80020";
		ram_buffer(4302) := X"88A90024";
		ram_buffer(4303) := X"88AA0028";
		ram_buffer(4304) := X"88AB002C";
		ram_buffer(4305) := X"88AC0030";
		ram_buffer(4306) := X"88AD0034";
		ram_buffer(4307) := X"88AE0038";
		ram_buffer(4308) := X"88AF003C";
		ram_buffer(4309) := X"98A80023";
		ram_buffer(4310) := X"98A90027";
		ram_buffer(4311) := X"98AA002B";
		ram_buffer(4312) := X"98AB002F";
		ram_buffer(4313) := X"98AC0033";
		ram_buffer(4314) := X"98AD0037";
		ram_buffer(4315) := X"98AE003B";
		ram_buffer(4316) := X"98AF003F";
		ram_buffer(4317) := X"AC880020";
		ram_buffer(4318) := X"AC890024";
		ram_buffer(4319) := X"AC8A0028";
		ram_buffer(4320) := X"AC8B002C";
		ram_buffer(4321) := X"AC8C0030";
		ram_buffer(4322) := X"AC8D0034";
		ram_buffer(4323) := X"AC8E0038";
		ram_buffer(4324) := X"AC8F003C";
		ram_buffer(4325) := X"24840040";
		ram_buffer(4326) := X"1487FFCE";
		ram_buffer(4327) := X"24A50040";
		ram_buffer(4328) := X"03003025";
		ram_buffer(4329) := X"30D8001F";
		ram_buffer(4330) := X"10D8001B";
		ram_buffer(4331) := X"00000000";
		ram_buffer(4332) := X"88A80000";
		ram_buffer(4333) := X"88A90004";
		ram_buffer(4334) := X"88AA0008";
		ram_buffer(4335) := X"88AB000C";
		ram_buffer(4336) := X"88AC0010";
		ram_buffer(4337) := X"88AD0014";
		ram_buffer(4338) := X"88AE0018";
		ram_buffer(4339) := X"88AF001C";
		ram_buffer(4340) := X"98A80003";
		ram_buffer(4341) := X"98A90007";
		ram_buffer(4342) := X"98AA000B";
		ram_buffer(4343) := X"98AB000F";
		ram_buffer(4344) := X"98AC0013";
		ram_buffer(4345) := X"98AD0017";
		ram_buffer(4346) := X"98AE001B";
		ram_buffer(4347) := X"98AF001F";
		ram_buffer(4348) := X"24A50020";
		ram_buffer(4349) := X"AC880000";
		ram_buffer(4350) := X"AC890004";
		ram_buffer(4351) := X"AC8A0008";
		ram_buffer(4352) := X"AC8B000C";
		ram_buffer(4353) := X"AC8C0010";
		ram_buffer(4354) := X"AC8D0014";
		ram_buffer(4355) := X"AC8E0018";
		ram_buffer(4356) := X"AC8F001C";
		ram_buffer(4357) := X"24840020";
		ram_buffer(4358) := X"33060003";
		ram_buffer(4359) := X"10D80008";
		ram_buffer(4360) := X"03063823";
		ram_buffer(4361) := X"00873821";
		ram_buffer(4362) := X"88A30000";
		ram_buffer(4363) := X"98A30003";
		ram_buffer(4364) := X"24840004";
		ram_buffer(4365) := X"24A50004";
		ram_buffer(4366) := X"1487FFFB";
		ram_buffer(4367) := X"AC83FFFC";
		ram_buffer(4368) := X"10C0FF87";
		ram_buffer(4369) := X"00863821";
		ram_buffer(4370) := X"80A30000";
		ram_buffer(4371) := X"24840001";
		ram_buffer(4372) := X"24A50001";
		ram_buffer(4373) := X"1487FFFC";
		ram_buffer(4374) := X"A083FFFF";
		ram_buffer(4375) := X"03E00008";
		ram_buffer(4376) := X"00000000";
		ram_buffer(4377) := X"28CA0008";
		ram_buffer(4378) := X"1540003E";
		ram_buffer(4379) := X"00801025";
		ram_buffer(4380) := X"10A00007";
		ram_buffer(4381) := X"00043823";
		ram_buffer(4382) := X"00000000";
		ram_buffer(4383) := X"30A500FF";
		ram_buffer(4384) := X"00055200";
		ram_buffer(4385) := X"00AA2825";
		ram_buffer(4386) := X"00055400";
		ram_buffer(4387) := X"00AA2825";
		ram_buffer(4388) := X"30EA0003";
		ram_buffer(4389) := X"11400003";
		ram_buffer(4390) := X"00CA3023";
		ram_buffer(4391) := X"A8850000";
		ram_buffer(4392) := X"008A2021";
		ram_buffer(4393) := X"30EA0004";
		ram_buffer(4394) := X"11400003";
		ram_buffer(4395) := X"00CA3023";
		ram_buffer(4396) := X"AC850000";
		ram_buffer(4397) := X"008A2021";
		ram_buffer(4398) := X"30D8003F";
		ram_buffer(4399) := X"10D80016";
		ram_buffer(4400) := X"00D83823";
		ram_buffer(4401) := X"00873821";
		ram_buffer(4402) := X"AC850000";
		ram_buffer(4403) := X"AC850004";
		ram_buffer(4404) := X"AC850008";
		ram_buffer(4405) := X"AC85000C";
		ram_buffer(4406) := X"AC850010";
		ram_buffer(4407) := X"AC850014";
		ram_buffer(4408) := X"AC850018";
		ram_buffer(4409) := X"AC85001C";
		ram_buffer(4410) := X"AC850020";
		ram_buffer(4411) := X"AC850024";
		ram_buffer(4412) := X"AC850028";
		ram_buffer(4413) := X"AC85002C";
		ram_buffer(4414) := X"AC850030";
		ram_buffer(4415) := X"AC850034";
		ram_buffer(4416) := X"AC850038";
		ram_buffer(4417) := X"AC85003C";
		ram_buffer(4418) := X"24840040";
		ram_buffer(4419) := X"1487FFEE";
		ram_buffer(4420) := X"00000000";
		ram_buffer(4421) := X"03003025";
		ram_buffer(4422) := X"30D8001F";
		ram_buffer(4423) := X"10D8000A";
		ram_buffer(4424) := X"00000000";
		ram_buffer(4425) := X"AC850000";
		ram_buffer(4426) := X"AC850004";
		ram_buffer(4427) := X"AC850008";
		ram_buffer(4428) := X"AC85000C";
		ram_buffer(4429) := X"AC850010";
		ram_buffer(4430) := X"AC850014";
		ram_buffer(4431) := X"AC850018";
		ram_buffer(4432) := X"AC85001C";
		ram_buffer(4433) := X"24840020";
		ram_buffer(4434) := X"33060003";
		ram_buffer(4435) := X"10D80005";
		ram_buffer(4436) := X"03063823";
		ram_buffer(4437) := X"00873821";
		ram_buffer(4438) := X"24840004";
		ram_buffer(4439) := X"1487FFFE";
		ram_buffer(4440) := X"AC85FFFC";
		ram_buffer(4441) := X"18C00004";
		ram_buffer(4442) := X"00863821";
		ram_buffer(4443) := X"24840001";
		ram_buffer(4444) := X"1487FFFE";
		ram_buffer(4445) := X"A085FFFF";
		ram_buffer(4446) := X"03E00008";
		ram_buffer(4447) := X"00000000";
		ram_buffer(4448) := X"24820001";
		ram_buffer(4449) := X"90830000";
		ram_buffer(4450) := X"00000000";
		ram_buffer(4451) := X"1460FFFD";
		ram_buffer(4452) := X"24840001";
		ram_buffer(4453) := X"03E00008";
		ram_buffer(4454) := X"00821023";
		ram_buffer(4455) := X"6D61696E";
		ram_buffer(4456) := X"00000000";
		ram_buffer(4457) := X"696E7075";
		ram_buffer(4458) := X"74000000";
		ram_buffer(4459) := X"74696D65";
		ram_buffer(4460) := X"00000000";
		ram_buffer(4461) := X"2E2E2F2E";
		ram_buffer(4462) := X"2E2F6672";
		ram_buffer(4463) := X"65657274";
		ram_buffer(4464) := X"6F732F71";
		ram_buffer(4465) := X"75657565";
		ram_buffer(4466) := X"2E630000";
		ram_buffer(4467) := X"2E2E2F2E";
		ram_buffer(4468) := X"2E2F6672";
		ram_buffer(4469) := X"65657274";
		ram_buffer(4470) := X"6F732F74";
		ram_buffer(4471) := X"61736B73";
		ram_buffer(4472) := X"2E630000";
		ram_buffer(4473) := X"49444C45";
		ram_buffer(4474) := X"00000000";
		ram_buffer(4475) := X"2E2E2F2E";
		ram_buffer(4476) := X"2E2F6672";
		ram_buffer(4477) := X"65657274";
		ram_buffer(4478) := X"6F732F70";
		ram_buffer(4479) := X"6F72742E";
		ram_buffer(4480) := X"63000000";
		ram_buffer(4481) := X"2E2E2F2E";
		ram_buffer(4482) := X"2E2F6672";
		ram_buffer(4483) := X"65657274";
		ram_buffer(4484) := X"6F732F68";
		ram_buffer(4485) := X"6561705F";
		ram_buffer(4486) := X"312E6300";
		ram_buffer(4487) := X"00000000";
		ram_buffer(4488) := X"00000000";
		ram_buffer(4489) := X"00000000";
		ram_buffer(4490) := X"00000000";
		ram_buffer(4491) := X"00000000";
		ram_buffer(4492) := X"00000000";
		ram_buffer(4493) := X"00000000";
		ram_buffer(4494) := X"00000000";
		ram_buffer(4495) := X"00000000";
		ram_buffer(4496) := X"00000000";
		ram_buffer(4497) := X"00000000";
		ram_buffer(4498) := X"00000000";
		ram_buffer(4499) := X"00000000";
		ram_buffer(4500) := X"00000000";
		ram_buffer(4501) := X"00000000";
		ram_buffer(4502) := X"00000000";
		ram_buffer(4503) := X"00000000";
		ram_buffer(4504) := X"00000000";
		ram_buffer(4505) := X"00000000";
		ram_buffer(4506) := X"00000000";
		ram_buffer(4507) := X"00000000";
		ram_buffer(4508) := X"00000000";
		ram_buffer(4509) := X"00000000";
		ram_buffer(4510) := X"00000000";
		ram_buffer(4511) := X"00000000";
		ram_buffer(4512) := X"00000000";
		ram_buffer(4513) := X"00000000";
		ram_buffer(4514) := X"00000000";
		ram_buffer(4515) := X"00000000";
		ram_buffer(4516) := X"00000000";
		ram_buffer(4517) := X"00000000";
		ram_buffer(4518) := X"00000000";
		ram_buffer(4519) := X"00000000";
		ram_buffer(4520) := X"00000000";
		ram_buffer(4521) := X"00000000";
		ram_buffer(4522) := X"00000000";
		ram_buffer(4523) := X"00000000";
		ram_buffer(4524) := X"00000000";
		ram_buffer(4525) := X"00000000";
		ram_buffer(4526) := X"00000000";
		ram_buffer(4527) := X"00000000";
		ram_buffer(4528) := X"00000000";
		ram_buffer(4529) := X"00000000";
		ram_buffer(4530) := X"00000000";
		ram_buffer(4531) := X"00000000";
		ram_buffer(4532) := X"00000000";
		ram_buffer(4533) := X"00000000";
		ram_buffer(4534) := X"00000000";
		ram_buffer(4535) := X"00000000";
		ram_buffer(4536) := X"00000000";
		ram_buffer(4537) := X"00000000";
		ram_buffer(4538) := X"00000000";
		ram_buffer(4539) := X"00000000";
		ram_buffer(4540) := X"00000000";
		ram_buffer(4541) := X"00000000";
		ram_buffer(4542) := X"00000000";
		ram_buffer(4543) := X"00000000";
		ram_buffer(4544) := X"00000000";
		ram_buffer(4545) := X"00000000";
		ram_buffer(4546) := X"00000000";
		ram_buffer(4547) := X"00000000";
		ram_buffer(4548) := X"00000000";
		ram_buffer(4549) := X"00000000";
		ram_buffer(4550) := X"00000000";
		ram_buffer(4551) := X"00000000";
		ram_buffer(4552) := X"00000000";
		ram_buffer(4553) := X"00000000";
		ram_buffer(4554) := X"00000000";
		ram_buffer(4555) := X"00000000";
		ram_buffer(4556) := X"00000000";
		ram_buffer(4557) := X"00000000";
		ram_buffer(4558) := X"00000000";
		ram_buffer(4559) := X"00000000";
		ram_buffer(4560) := X"00000000";
		ram_buffer(4561) := X"00000000";
		ram_buffer(4562) := X"00000000";
		ram_buffer(4563) := X"00000000";
		ram_buffer(4564) := X"00000000";
		ram_buffer(4565) := X"00000000";
		ram_buffer(4566) := X"00000000";
		ram_buffer(4567) := X"00000000";
		ram_buffer(4568) := X"00000000";
		ram_buffer(4569) := X"00000000";
		ram_buffer(4570) := X"00000000";
		ram_buffer(4571) := X"00000000";
		ram_buffer(4572) := X"00000000";
		ram_buffer(4573) := X"00000000";
		ram_buffer(4574) := X"00000000";
		ram_buffer(4575) := X"00000000";
		ram_buffer(4576) := X"00000000";
		ram_buffer(4577) := X"00000000";
		ram_buffer(4578) := X"00000000";
		ram_buffer(4579) := X"00000000";
		ram_buffer(4580) := X"00000000";
		ram_buffer(4581) := X"00000000";
		ram_buffer(4582) := X"00000000";
		ram_buffer(4583) := X"00000000";
		ram_buffer(4584) := X"00000000";
		ram_buffer(4585) := X"00000000";
		ram_buffer(4586) := X"00000000";
		ram_buffer(4587) := X"00000000";
		ram_buffer(4588) := X"00000000";
		ram_buffer(4589) := X"00000000";
		ram_buffer(4590) := X"00000000";
		ram_buffer(4591) := X"00000000";
		ram_buffer(4592) := X"00000000";
		ram_buffer(4593) := X"00000000";
		ram_buffer(4594) := X"00000000";
		ram_buffer(4595) := X"00000000";
		ram_buffer(4596) := X"00000000";
		ram_buffer(4597) := X"00000000";
		ram_buffer(4598) := X"00000000";
		ram_buffer(4599) := X"00000000";
		ram_buffer(4600) := X"00000000";
		ram_buffer(4601) := X"00000000";
		ram_buffer(4602) := X"00000000";
		ram_buffer(4603) := X"00000000";
		ram_buffer(4604) := X"00000000";
		ram_buffer(4605) := X"00000000";
		ram_buffer(4606) := X"00000000";
		ram_buffer(4607) := X"00000000";
		ram_buffer(4608) := X"00000000";
		ram_buffer(4609) := X"00000000";
		ram_buffer(4610) := X"00000000";
		ram_buffer(4611) := X"00000000";
		ram_buffer(4612) := X"00000000";
		ram_buffer(4613) := X"00000000";
		ram_buffer(4614) := X"00000000";
		ram_buffer(4615) := X"00000000";
		ram_buffer(4616) := X"00000000";
		ram_buffer(4617) := X"00000000";
		ram_buffer(4618) := X"00000000";
		ram_buffer(4619) := X"00000000";
		ram_buffer(4620) := X"00000000";
		ram_buffer(4621) := X"00000000";
		ram_buffer(4622) := X"00000000";
		ram_buffer(4623) := X"00000000";
		ram_buffer(4624) := X"00000000";
		ram_buffer(4625) := X"00000000";
		ram_buffer(4626) := X"00000000";
		ram_buffer(4627) := X"00000000";
		ram_buffer(4628) := X"00000000";
		ram_buffer(4629) := X"00000000";
		ram_buffer(4630) := X"00000000";
		ram_buffer(4631) := X"00000000";
		ram_buffer(4632) := X"00000000";
		ram_buffer(4633) := X"00000000";
		ram_buffer(4634) := X"00000000";
		ram_buffer(4635) := X"00000000";
		ram_buffer(4636) := X"00000000";
		ram_buffer(4637) := X"00000000";
		ram_buffer(4638) := X"00000000";
		ram_buffer(4639) := X"00000000";
		ram_buffer(4640) := X"00000000";
		ram_buffer(4641) := X"00000000";
		ram_buffer(4642) := X"00000000";
		ram_buffer(4643) := X"00000000";
		ram_buffer(4644) := X"00000000";
		ram_buffer(4645) := X"00000000";
		ram_buffer(4646) := X"00000000";
		ram_buffer(4647) := X"00000000";
		ram_buffer(4648) := X"00000000";
		ram_buffer(4649) := X"00000000";
		ram_buffer(4650) := X"00000000";
		ram_buffer(4651) := X"00000000";
		ram_buffer(4652) := X"00000000";
		ram_buffer(4653) := X"00000000";
		ram_buffer(4654) := X"00000000";
		ram_buffer(4655) := X"00000000";
		ram_buffer(4656) := X"00000000";
		ram_buffer(4657) := X"00000000";
		ram_buffer(4658) := X"00000000";
		ram_buffer(4659) := X"00000000";
		ram_buffer(4660) := X"00000000";
		ram_buffer(4661) := X"00000000";
		ram_buffer(4662) := X"00000000";
		ram_buffer(4663) := X"00000000";
		ram_buffer(4664) := X"00000000";
		ram_buffer(4665) := X"00000000";
		ram_buffer(4666) := X"00000000";
		ram_buffer(4667) := X"00000000";
		ram_buffer(4668) := X"00000000";
		ram_buffer(4669) := X"00000000";
		ram_buffer(4670) := X"00000000";
		ram_buffer(4671) := X"00000000";
		ram_buffer(4672) := X"00000000";
		ram_buffer(4673) := X"00000000";
		ram_buffer(4674) := X"00000000";
		ram_buffer(4675) := X"00000000";
		ram_buffer(4676) := X"00000000";
		ram_buffer(4677) := X"00000000";
		ram_buffer(4678) := X"00000000";
		ram_buffer(4679) := X"00000000";
		ram_buffer(4680) := X"00000000";
		ram_buffer(4681) := X"00000000";
		ram_buffer(4682) := X"00000000";
		ram_buffer(4683) := X"00000000";
		ram_buffer(4684) := X"00000000";
		ram_buffer(4685) := X"00000000";
		ram_buffer(4686) := X"00000000";
		ram_buffer(4687) := X"00000000";
		ram_buffer(4688) := X"00000000";
		ram_buffer(4689) := X"00000000";
		ram_buffer(4690) := X"00000000";
		ram_buffer(4691) := X"00000000";
		ram_buffer(4692) := X"00000000";
		ram_buffer(4693) := X"00000000";
		ram_buffer(4694) := X"00000000";
		ram_buffer(4695) := X"00000000";
		ram_buffer(4696) := X"00000000";
		ram_buffer(4697) := X"00000000";
		ram_buffer(4698) := X"00000000";
		ram_buffer(4699) := X"00000000";
		ram_buffer(4700) := X"00000000";
		ram_buffer(4701) := X"00000000";
		ram_buffer(4702) := X"00000000";
		ram_buffer(4703) := X"00000000";
		ram_buffer(4704) := X"00000000";
		ram_buffer(4705) := X"00000000";
		ram_buffer(4706) := X"00000000";
		ram_buffer(4707) := X"00000000";
		ram_buffer(4708) := X"00000000";
		ram_buffer(4709) := X"00000000";
		ram_buffer(4710) := X"00000000";
		ram_buffer(4711) := X"00000000";
		ram_buffer(4712) := X"00000000";
		ram_buffer(4713) := X"00000000";
		ram_buffer(4714) := X"00000000";
		ram_buffer(4715) := X"00000000";
		ram_buffer(4716) := X"00000000";
		ram_buffer(4717) := X"00000000";
		ram_buffer(4718) := X"00000000";
		ram_buffer(4719) := X"00000000";
		ram_buffer(4720) := X"00000000";
		ram_buffer(4721) := X"00000000";
		ram_buffer(4722) := X"00000000";
		ram_buffer(4723) := X"00000000";
		ram_buffer(4724) := X"00000000";
		ram_buffer(4725) := X"00000000";
		ram_buffer(4726) := X"00000000";
		ram_buffer(4727) := X"00000000";
		ram_buffer(4728) := X"00000000";
		ram_buffer(4729) := X"00000000";
		ram_buffer(4730) := X"00000000";
		ram_buffer(4731) := X"00000000";
		ram_buffer(4732) := X"00000000";
		ram_buffer(4733) := X"00000000";
		ram_buffer(4734) := X"00000000";
		ram_buffer(4735) := X"00000000";
		ram_buffer(4736) := X"00000000";
		ram_buffer(4737) := X"00000000";
		ram_buffer(4738) := X"00000000";
		ram_buffer(4739) := X"00000000";
		ram_buffer(4740) := X"00000000";
		ram_buffer(4741) := X"00000000";
		ram_buffer(4742) := X"00000000";
		ram_buffer(4743) := X"00000000";
		ram_buffer(4744) := X"00000000";
		ram_buffer(4745) := X"00000000";
		ram_buffer(4746) := X"00000000";
		ram_buffer(4747) := X"00000000";
		ram_buffer(4748) := X"00000000";
		ram_buffer(4749) := X"00000000";
		ram_buffer(4750) := X"00000000";
		ram_buffer(4751) := X"00000000";
		ram_buffer(4752) := X"00000000";
		ram_buffer(4753) := X"00000000";
		ram_buffer(4754) := X"00000000";
		ram_buffer(4755) := X"00000000";
		ram_buffer(4756) := X"00000000";
		ram_buffer(4757) := X"00000000";
		ram_buffer(4758) := X"00000000";
		ram_buffer(4759) := X"00000000";
		ram_buffer(4760) := X"00000000";
		ram_buffer(4761) := X"00000000";
		ram_buffer(4762) := X"00000000";
		ram_buffer(4763) := X"00000000";
		ram_buffer(4764) := X"00000000";
		ram_buffer(4765) := X"00000000";
		ram_buffer(4766) := X"00000000";
		ram_buffer(4767) := X"00000000";
		ram_buffer(4768) := X"00000000";
		ram_buffer(4769) := X"00000000";
		ram_buffer(4770) := X"00000000";
		ram_buffer(4771) := X"00000000";
		ram_buffer(4772) := X"00000000";
		ram_buffer(4773) := X"00000000";
		ram_buffer(4774) := X"00000000";
		ram_buffer(4775) := X"00000000";
		ram_buffer(4776) := X"00000000";
		ram_buffer(4777) := X"00000000";
		ram_buffer(4778) := X"00000000";
		ram_buffer(4779) := X"00000000";
		ram_buffer(4780) := X"00000000";
		ram_buffer(4781) := X"00000000";
		ram_buffer(4782) := X"00000000";
		ram_buffer(4783) := X"00000000";
		ram_buffer(4784) := X"00000000";
		ram_buffer(4785) := X"00000000";
		ram_buffer(4786) := X"00000000";
		ram_buffer(4787) := X"00000000";
		ram_buffer(4788) := X"00000000";
		ram_buffer(4789) := X"00000000";
		ram_buffer(4790) := X"00000000";
		ram_buffer(4791) := X"00000000";
		ram_buffer(4792) := X"00000000";
		ram_buffer(4793) := X"00000000";
		ram_buffer(4794) := X"00000000";
		ram_buffer(4795) := X"00000000";
		ram_buffer(4796) := X"00000000";
		ram_buffer(4797) := X"00000000";
		ram_buffer(4798) := X"00000000";
		ram_buffer(4799) := X"00000000";
		ram_buffer(4800) := X"00000000";
		ram_buffer(4801) := X"00000000";
		ram_buffer(4802) := X"00000000";
		ram_buffer(4803) := X"00000000";
		ram_buffer(4804) := X"00000000";
		ram_buffer(4805) := X"00000000";
		ram_buffer(4806) := X"00000000";
		ram_buffer(4807) := X"00000000";
		ram_buffer(4808) := X"00000000";
		ram_buffer(4809) := X"00000000";
		ram_buffer(4810) := X"00000000";
		ram_buffer(4811) := X"00000000";
		ram_buffer(4812) := X"00000000";
		ram_buffer(4813) := X"00000000";
		ram_buffer(4814) := X"00000000";
		ram_buffer(4815) := X"00000000";
		ram_buffer(4816) := X"00000000";
		ram_buffer(4817) := X"00000000";
		ram_buffer(4818) := X"00000000";
		ram_buffer(4819) := X"00000000";
		ram_buffer(4820) := X"00000000";
		ram_buffer(4821) := X"00000000";
		ram_buffer(4822) := X"00000000";
		ram_buffer(4823) := X"00000000";
		ram_buffer(4824) := X"00000000";
		ram_buffer(4825) := X"00000000";
		ram_buffer(4826) := X"00000000";
		ram_buffer(4827) := X"00000000";
		ram_buffer(4828) := X"00000000";
		ram_buffer(4829) := X"00000000";
		ram_buffer(4830) := X"00000000";
		ram_buffer(4831) := X"00000000";
		ram_buffer(4832) := X"00000000";
		ram_buffer(4833) := X"00000000";
		ram_buffer(4834) := X"00000000";
		ram_buffer(4835) := X"00000000";
		ram_buffer(4836) := X"00000000";
		ram_buffer(4837) := X"00000000";
		ram_buffer(4838) := X"00000000";
		ram_buffer(4839) := X"00000000";
		ram_buffer(4840) := X"00000000";
		ram_buffer(4841) := X"00000000";
		ram_buffer(4842) := X"00000000";
		ram_buffer(4843) := X"00000000";
		ram_buffer(4844) := X"00000000";
		ram_buffer(4845) := X"00000000";
		ram_buffer(4846) := X"00000000";
		ram_buffer(4847) := X"00000000";
		ram_buffer(4848) := X"00000000";
		ram_buffer(4849) := X"00000000";
		ram_buffer(4850) := X"00000000";
		ram_buffer(4851) := X"00000000";
		ram_buffer(4852) := X"00000000";
		ram_buffer(4853) := X"00000000";
		ram_buffer(4854) := X"00000000";
		ram_buffer(4855) := X"00000000";
		ram_buffer(4856) := X"00000000";
		ram_buffer(4857) := X"00000000";
		ram_buffer(4858) := X"00000000";
		ram_buffer(4859) := X"00000000";
		ram_buffer(4860) := X"00000000";
		ram_buffer(4861) := X"00000000";
		ram_buffer(4862) := X"00000000";
		ram_buffer(4863) := X"00000000";
		ram_buffer(4864) := X"00000000";
		ram_buffer(4865) := X"00000000";
		ram_buffer(4866) := X"00000000";
		ram_buffer(4867) := X"00000000";
		ram_buffer(4868) := X"00000000";
		ram_buffer(4869) := X"00000000";
		ram_buffer(4870) := X"00000000";
		ram_buffer(4871) := X"00000000";
		ram_buffer(4872) := X"00000000";
		ram_buffer(4873) := X"00000000";
		ram_buffer(4874) := X"00000000";
		ram_buffer(4875) := X"00000000";
		ram_buffer(4876) := X"00000000";
		ram_buffer(4877) := X"00000000";
		ram_buffer(4878) := X"00000000";
		ram_buffer(4879) := X"00000000";
		ram_buffer(4880) := X"00000000";
		ram_buffer(4881) := X"00000000";
		ram_buffer(4882) := X"00000000";
		ram_buffer(4883) := X"00000000";
		ram_buffer(4884) := X"00000000";
		ram_buffer(4885) := X"00000000";
		ram_buffer(4886) := X"00000000";
		ram_buffer(4887) := X"00000000";
		ram_buffer(4888) := X"00000000";
		ram_buffer(4889) := X"00000000";
		ram_buffer(4890) := X"00000000";
		ram_buffer(4891) := X"00000000";
		ram_buffer(4892) := X"00000000";
		ram_buffer(4893) := X"00000000";
		ram_buffer(4894) := X"00000000";
		ram_buffer(4895) := X"00000000";
		ram_buffer(4896) := X"00000000";
		ram_buffer(4897) := X"00000000";
		ram_buffer(4898) := X"00000000";
		ram_buffer(4899) := X"00000000";
		ram_buffer(4900) := X"00000000";
		ram_buffer(4901) := X"00000000";
		ram_buffer(4902) := X"00000000";
		ram_buffer(4903) := X"00000000";
		ram_buffer(4904) := X"00000000";
		ram_buffer(4905) := X"00000000";
		ram_buffer(4906) := X"00000000";
		ram_buffer(4907) := X"00000000";
		ram_buffer(4908) := X"00000000";
		ram_buffer(4909) := X"00000000";
		ram_buffer(4910) := X"00000000";
		ram_buffer(4911) := X"00000000";
		ram_buffer(4912) := X"00000000";
		ram_buffer(4913) := X"00000000";
		ram_buffer(4914) := X"00000000";
		ram_buffer(4915) := X"00000000";
		ram_buffer(4916) := X"00000000";
		ram_buffer(4917) := X"00000000";
		ram_buffer(4918) := X"00000000";
		ram_buffer(4919) := X"00000000";
		ram_buffer(4920) := X"00000000";
		ram_buffer(4921) := X"00000000";
		ram_buffer(4922) := X"00000000";
		ram_buffer(4923) := X"00000000";
		ram_buffer(4924) := X"00000000";
		ram_buffer(4925) := X"00000000";
		ram_buffer(4926) := X"00000000";
		ram_buffer(4927) := X"00000000";
		ram_buffer(4928) := X"00000000";
		ram_buffer(4929) := X"00000000";
		ram_buffer(4930) := X"00000000";
		ram_buffer(4931) := X"00000000";
		ram_buffer(4932) := X"00000000";
		ram_buffer(4933) := X"00000000";
		ram_buffer(4934) := X"00000000";
		ram_buffer(4935) := X"00000000";
		ram_buffer(4936) := X"00000000";
		ram_buffer(4937) := X"00000000";
		ram_buffer(4938) := X"00000000";
		ram_buffer(4939) := X"00000000";
		ram_buffer(4940) := X"00000000";
		ram_buffer(4941) := X"00000000";
		ram_buffer(4942) := X"00000000";
		ram_buffer(4943) := X"00000000";
		ram_buffer(4944) := X"00000000";
		ram_buffer(4945) := X"00000000";
		ram_buffer(4946) := X"00000000";
		ram_buffer(4947) := X"00000000";
		ram_buffer(4948) := X"00000000";
		ram_buffer(4949) := X"00000000";
		ram_buffer(4950) := X"00000000";
		ram_buffer(4951) := X"00000000";
		ram_buffer(4952) := X"00000000";
		ram_buffer(4953) := X"00000000";
		ram_buffer(4954) := X"00000000";
		ram_buffer(4955) := X"00000000";
		ram_buffer(4956) := X"00000000";
		ram_buffer(4957) := X"00000000";
		ram_buffer(4958) := X"00000000";
		ram_buffer(4959) := X"00000000";
		ram_buffer(4960) := X"00000000";
		ram_buffer(4961) := X"00000000";
		ram_buffer(4962) := X"00000000";
		ram_buffer(4963) := X"00000000";
		ram_buffer(4964) := X"00000000";
		ram_buffer(4965) := X"00000000";
		ram_buffer(4966) := X"00000000";
		ram_buffer(4967) := X"00000000";
		ram_buffer(4968) := X"00000000";
		ram_buffer(4969) := X"00000000";
		ram_buffer(4970) := X"00000000";
		ram_buffer(4971) := X"00000000";
		ram_buffer(4972) := X"00000000";
		ram_buffer(4973) := X"00000000";
		ram_buffer(4974) := X"00000000";
		ram_buffer(4975) := X"00000000";
		ram_buffer(4976) := X"00000000";
		ram_buffer(4977) := X"00000000";
		ram_buffer(4978) := X"00000000";
		ram_buffer(4979) := X"00000000";
		ram_buffer(4980) := X"00000000";
		ram_buffer(4981) := X"00000000";
		ram_buffer(4982) := X"00000000";
		ram_buffer(4983) := X"00000000";
		ram_buffer(4984) := X"00000000";
		ram_buffer(4985) := X"00000000";
		ram_buffer(4986) := X"00000000";
		ram_buffer(4987) := X"00000000";
		ram_buffer(4988) := X"00000000";
		ram_buffer(4989) := X"00000000";
		ram_buffer(4990) := X"00000000";
		ram_buffer(4991) := X"00000000";
		ram_buffer(4992) := X"00000000";
		ram_buffer(4993) := X"00000000";
		ram_buffer(4994) := X"00000000";
		ram_buffer(4995) := X"00000000";
		ram_buffer(4996) := X"00000000";
		ram_buffer(4997) := X"00000000";
		ram_buffer(4998) := X"00000000";
		ram_buffer(4999) := X"00000000";
		ram_buffer(5000) := X"00000000";
		ram_buffer(5001) := X"00000000";
		ram_buffer(5002) := X"00000000";
		ram_buffer(5003) := X"00000000";
		ram_buffer(5004) := X"00000000";
		ram_buffer(5005) := X"00000000";
		ram_buffer(5006) := X"00000000";
		ram_buffer(5007) := X"00000000";
		ram_buffer(5008) := X"00000000";
		ram_buffer(5009) := X"00000000";
		ram_buffer(5010) := X"00000000";
		ram_buffer(5011) := X"00000000";
		ram_buffer(5012) := X"00000000";
		ram_buffer(5013) := X"00000000";
		ram_buffer(5014) := X"00000000";
		ram_buffer(5015) := X"00000000";
		ram_buffer(5016) := X"00000000";
		ram_buffer(5017) := X"00000000";
		ram_buffer(5018) := X"00000000";
		ram_buffer(5019) := X"00000000";
		ram_buffer(5020) := X"00000000";
		ram_buffer(5021) := X"00000000";
		ram_buffer(5022) := X"00000000";
		ram_buffer(5023) := X"00000000";
		ram_buffer(5024) := X"00000000";
		ram_buffer(5025) := X"00000000";
		ram_buffer(5026) := X"00000000";
		ram_buffer(5027) := X"00000000";
		ram_buffer(5028) := X"00000000";
		ram_buffer(5029) := X"00000000";
		ram_buffer(5030) := X"00000000";
		ram_buffer(5031) := X"00000000";
		ram_buffer(5032) := X"00000000";
		ram_buffer(5033) := X"00000000";
		ram_buffer(5034) := X"00000000";
		ram_buffer(5035) := X"00000000";
		ram_buffer(5036) := X"00000000";
		ram_buffer(5037) := X"00000000";
		ram_buffer(5038) := X"00000000";
		ram_buffer(5039) := X"00000000";
		ram_buffer(5040) := X"00000000";
		ram_buffer(5041) := X"00000000";
		ram_buffer(5042) := X"00000000";
		ram_buffer(5043) := X"00000000";
		ram_buffer(5044) := X"00000000";
		ram_buffer(5045) := X"00000000";
		ram_buffer(5046) := X"00000000";
		ram_buffer(5047) := X"00000000";
		ram_buffer(5048) := X"00000000";
		ram_buffer(5049) := X"00000000";
		ram_buffer(5050) := X"00000000";
		ram_buffer(5051) := X"00000000";
		ram_buffer(5052) := X"00000000";
		ram_buffer(5053) := X"00000000";
		ram_buffer(5054) := X"00000000";
		ram_buffer(5055) := X"00000000";
		ram_buffer(5056) := X"00000000";
		ram_buffer(5057) := X"00000000";
		ram_buffer(5058) := X"00000000";
		ram_buffer(5059) := X"00000000";
		ram_buffer(5060) := X"00000000";
		ram_buffer(5061) := X"00000000";
		ram_buffer(5062) := X"00000000";
		ram_buffer(5063) := X"00000000";
		ram_buffer(5064) := X"00000000";
		ram_buffer(5065) := X"00000000";
		ram_buffer(5066) := X"00000000";
		ram_buffer(5067) := X"00000000";
		ram_buffer(5068) := X"00000000";
		ram_buffer(5069) := X"00000000";
		ram_buffer(5070) := X"00000000";
		ram_buffer(5071) := X"00000000";
		ram_buffer(5072) := X"00000000";
		ram_buffer(5073) := X"00000000";
		ram_buffer(5074) := X"00000000";
		ram_buffer(5075) := X"00000000";
		ram_buffer(5076) := X"00000000";
		ram_buffer(5077) := X"00000000";
		ram_buffer(5078) := X"00000000";
		ram_buffer(5079) := X"00000000";
		ram_buffer(5080) := X"00000000";
		ram_buffer(5081) := X"00000000";
		ram_buffer(5082) := X"00000000";
		ram_buffer(5083) := X"00000000";
		ram_buffer(5084) := X"00000000";
		ram_buffer(5085) := X"00000000";
		ram_buffer(5086) := X"00000000";
		ram_buffer(5087) := X"00000000";
		ram_buffer(5088) := X"00000000";
		ram_buffer(5089) := X"00000000";
		ram_buffer(5090) := X"00000000";
		ram_buffer(5091) := X"00000000";
		ram_buffer(5092) := X"00000000";
		ram_buffer(5093) := X"00000000";
		ram_buffer(5094) := X"00000000";
		ram_buffer(5095) := X"00000000";
		ram_buffer(5096) := X"00000000";
		ram_buffer(5097) := X"00000000";
		ram_buffer(5098) := X"00000000";
		ram_buffer(5099) := X"00000000";
		ram_buffer(5100) := X"00000000";
		ram_buffer(5101) := X"00000000";
		ram_buffer(5102) := X"00000000";
		ram_buffer(5103) := X"00000000";
		ram_buffer(5104) := X"00000000";
		ram_buffer(5105) := X"00000000";
		ram_buffer(5106) := X"00000000";
		ram_buffer(5107) := X"00000000";
		ram_buffer(5108) := X"00000000";
		ram_buffer(5109) := X"00000000";
		ram_buffer(5110) := X"00000000";
		ram_buffer(5111) := X"00000000";
		ram_buffer(5112) := X"00000000";
		ram_buffer(5113) := X"00000000";
		ram_buffer(5114) := X"00000000";
		ram_buffer(5115) := X"00000000";
		ram_buffer(5116) := X"00000000";
		ram_buffer(5117) := X"00000000";
		ram_buffer(5118) := X"00000000";
		ram_buffer(5119) := X"00000000";
		ram_buffer(5120) := X"00000000";
		ram_buffer(5121) := X"00000000";
		ram_buffer(5122) := X"00000000";
		ram_buffer(5123) := X"00000000";
		ram_buffer(5124) := X"00000000";
		ram_buffer(5125) := X"00000000";
		ram_buffer(5126) := X"00000000";
		ram_buffer(5127) := X"00000000";
		ram_buffer(5128) := X"00000000";
		ram_buffer(5129) := X"00000000";
		ram_buffer(5130) := X"00000000";
		ram_buffer(5131) := X"00000000";
		ram_buffer(5132) := X"00000000";
		ram_buffer(5133) := X"00000000";
		ram_buffer(5134) := X"00000000";
		ram_buffer(5135) := X"00000000";
		ram_buffer(5136) := X"00000000";
		ram_buffer(5137) := X"00000000";
		ram_buffer(5138) := X"00000000";
		ram_buffer(5139) := X"00000000";
		ram_buffer(5140) := X"00000000";
		ram_buffer(5141) := X"00000000";
		ram_buffer(5142) := X"00000000";
		ram_buffer(5143) := X"00000000";
		ram_buffer(5144) := X"00000000";
		ram_buffer(5145) := X"00000000";
		ram_buffer(5146) := X"00000000";
		ram_buffer(5147) := X"00000000";
		ram_buffer(5148) := X"00000000";
		ram_buffer(5149) := X"00000000";
		ram_buffer(5150) := X"00000000";
		ram_buffer(5151) := X"00000000";
		ram_buffer(5152) := X"00000000";
		ram_buffer(5153) := X"00000000";
		ram_buffer(5154) := X"00000000";
		ram_buffer(5155) := X"00000000";
		ram_buffer(5156) := X"00000000";
		ram_buffer(5157) := X"00000000";
		ram_buffer(5158) := X"00000000";
		ram_buffer(5159) := X"00000000";
		ram_buffer(5160) := X"00000000";
		ram_buffer(5161) := X"00000000";
		ram_buffer(5162) := X"00000000";
		ram_buffer(5163) := X"00000000";
		ram_buffer(5164) := X"00000000";
		ram_buffer(5165) := X"00000000";
		ram_buffer(5166) := X"00000000";
		ram_buffer(5167) := X"00000000";
		ram_buffer(5168) := X"00000000";
		ram_buffer(5169) := X"00000000";
		ram_buffer(5170) := X"00000000";
		ram_buffer(5171) := X"00000000";
		ram_buffer(5172) := X"00000000";
		ram_buffer(5173) := X"00000000";
		ram_buffer(5174) := X"00000000";
		ram_buffer(5175) := X"00000000";
		ram_buffer(5176) := X"00000000";
		ram_buffer(5177) := X"00000000";
		ram_buffer(5178) := X"00000000";
		ram_buffer(5179) := X"00000000";
		ram_buffer(5180) := X"00000000";
		ram_buffer(5181) := X"00000000";
		ram_buffer(5182) := X"00000000";
		ram_buffer(5183) := X"00000000";
		ram_buffer(5184) := X"00000000";
		ram_buffer(5185) := X"00000000";
		ram_buffer(5186) := X"00000000";
		ram_buffer(5187) := X"00000000";
		ram_buffer(5188) := X"00000000";
		ram_buffer(5189) := X"00000000";
		ram_buffer(5190) := X"00000000";
		ram_buffer(5191) := X"00000000";
		ram_buffer(5192) := X"00000000";
		ram_buffer(5193) := X"00000000";
		ram_buffer(5194) := X"00000000";
		ram_buffer(5195) := X"00000000";
		ram_buffer(5196) := X"00000000";
		ram_buffer(5197) := X"00000000";
		ram_buffer(5198) := X"00000000";
		ram_buffer(5199) := X"00000000";
		ram_buffer(5200) := X"00000000";
		ram_buffer(5201) := X"00000000";
		ram_buffer(5202) := X"00000000";
		ram_buffer(5203) := X"00000000";
		ram_buffer(5204) := X"00000000";
		ram_buffer(5205) := X"00000000";
		ram_buffer(5206) := X"00000000";
		ram_buffer(5207) := X"00000000";
		ram_buffer(5208) := X"00000000";
		ram_buffer(5209) := X"00000000";
		ram_buffer(5210) := X"00000000";
		ram_buffer(5211) := X"00000000";
		ram_buffer(5212) := X"00000000";
		ram_buffer(5213) := X"00000000";
		ram_buffer(5214) := X"00000000";
		ram_buffer(5215) := X"00000000";
		ram_buffer(5216) := X"00000000";
		ram_buffer(5217) := X"00000000";
		ram_buffer(5218) := X"00000000";
		ram_buffer(5219) := X"00000000";
		ram_buffer(5220) := X"00000000";
		ram_buffer(5221) := X"00000000";
		ram_buffer(5222) := X"00000000";
		ram_buffer(5223) := X"00000000";
		ram_buffer(5224) := X"00000000";
		ram_buffer(5225) := X"00000000";
		ram_buffer(5226) := X"00000000";
		ram_buffer(5227) := X"00000000";
		ram_buffer(5228) := X"00000000";
		ram_buffer(5229) := X"00000000";
		ram_buffer(5230) := X"00000000";
		ram_buffer(5231) := X"00000000";
		ram_buffer(5232) := X"00000000";
		ram_buffer(5233) := X"00000000";
		ram_buffer(5234) := X"00000000";
		ram_buffer(5235) := X"00000000";
		ram_buffer(5236) := X"00000000";
		ram_buffer(5237) := X"00000000";
		ram_buffer(5238) := X"00000000";
		ram_buffer(5239) := X"00000000";
		ram_buffer(5240) := X"00000000";
		ram_buffer(5241) := X"00000000";
		ram_buffer(5242) := X"00000000";
		ram_buffer(5243) := X"00000000";
		ram_buffer(5244) := X"00000000";
		ram_buffer(5245) := X"00000000";
		ram_buffer(5246) := X"00000000";
		ram_buffer(5247) := X"00000000";
		ram_buffer(5248) := X"00000000";
		ram_buffer(5249) := X"00000000";
		ram_buffer(5250) := X"00000000";
		ram_buffer(5251) := X"00000000";
		ram_buffer(5252) := X"00000000";
		ram_buffer(5253) := X"00000000";
		ram_buffer(5254) := X"00000000";
		ram_buffer(5255) := X"00000000";
		ram_buffer(5256) := X"00000000";
		ram_buffer(5257) := X"00000000";
		ram_buffer(5258) := X"00000000";
		ram_buffer(5259) := X"00000000";
		ram_buffer(5260) := X"00000000";
		ram_buffer(5261) := X"00000000";
		ram_buffer(5262) := X"00000000";
		ram_buffer(5263) := X"00000000";
		ram_buffer(5264) := X"00000000";
		ram_buffer(5265) := X"00000000";
		ram_buffer(5266) := X"00000000";
		ram_buffer(5267) := X"00000000";
		ram_buffer(5268) := X"00000000";
		ram_buffer(5269) := X"00000000";
		ram_buffer(5270) := X"00000000";
		ram_buffer(5271) := X"00000000";
		ram_buffer(5272) := X"00000000";
		ram_buffer(5273) := X"00000000";
		ram_buffer(5274) := X"00000000";
		ram_buffer(5275) := X"00000000";
		ram_buffer(5276) := X"00000000";
		ram_buffer(5277) := X"00000000";
		ram_buffer(5278) := X"00000000";
		ram_buffer(5279) := X"00000000";
		ram_buffer(5280) := X"00000000";
		ram_buffer(5281) := X"00000000";
		ram_buffer(5282) := X"00000000";
		ram_buffer(5283) := X"00000000";
		ram_buffer(5284) := X"00000000";
		ram_buffer(5285) := X"00000000";
		ram_buffer(5286) := X"00000000";
		ram_buffer(5287) := X"00000000";
		ram_buffer(5288) := X"00000000";
		ram_buffer(5289) := X"00000000";
		ram_buffer(5290) := X"00000000";
		ram_buffer(5291) := X"00000000";
		ram_buffer(5292) := X"00000000";
		ram_buffer(5293) := X"00000000";
		ram_buffer(5294) := X"00000000";
		ram_buffer(5295) := X"00000000";
		ram_buffer(5296) := X"00000000";
		ram_buffer(5297) := X"00000000";
		ram_buffer(5298) := X"00000000";
		ram_buffer(5299) := X"00000000";
		ram_buffer(5300) := X"00000000";
		ram_buffer(5301) := X"00000000";
		ram_buffer(5302) := X"00000000";
		ram_buffer(5303) := X"00000000";
		ram_buffer(5304) := X"00000000";
		ram_buffer(5305) := X"00000000";
		ram_buffer(5306) := X"00000000";
		ram_buffer(5307) := X"00000000";
		ram_buffer(5308) := X"00000000";
		ram_buffer(5309) := X"00000000";
		ram_buffer(5310) := X"00000000";
		ram_buffer(5311) := X"00000000";
		ram_buffer(5312) := X"00000000";
		ram_buffer(5313) := X"00000000";
		ram_buffer(5314) := X"00000000";
		ram_buffer(5315) := X"00000000";
		ram_buffer(5316) := X"00000000";
		ram_buffer(5317) := X"00000000";
		ram_buffer(5318) := X"00000000";
		ram_buffer(5319) := X"00000000";
		ram_buffer(5320) := X"00000000";
		ram_buffer(5321) := X"00000000";
		ram_buffer(5322) := X"00000000";
		ram_buffer(5323) := X"00000000";
		ram_buffer(5324) := X"00000000";
		ram_buffer(5325) := X"00000000";
		ram_buffer(5326) := X"00000000";
		ram_buffer(5327) := X"00000000";
		ram_buffer(5328) := X"00000000";
		ram_buffer(5329) := X"00000000";
		ram_buffer(5330) := X"00000000";
		ram_buffer(5331) := X"00000000";
		ram_buffer(5332) := X"00000000";
		ram_buffer(5333) := X"00000000";
		ram_buffer(5334) := X"00000000";
		ram_buffer(5335) := X"00000000";
		ram_buffer(5336) := X"00000000";
		ram_buffer(5337) := X"00000000";
		ram_buffer(5338) := X"00000000";
		ram_buffer(5339) := X"00000000";
		ram_buffer(5340) := X"00000000";
		ram_buffer(5341) := X"00000000";
		ram_buffer(5342) := X"00000000";
		ram_buffer(5343) := X"00000000";
		ram_buffer(5344) := X"00000000";
		ram_buffer(5345) := X"00000000";
		ram_buffer(5346) := X"00000000";
		ram_buffer(5347) := X"00000000";
		ram_buffer(5348) := X"00000000";
		ram_buffer(5349) := X"00000000";
		ram_buffer(5350) := X"00000000";
		ram_buffer(5351) := X"00000000";
		ram_buffer(5352) := X"00000000";
		ram_buffer(5353) := X"00000000";
		ram_buffer(5354) := X"00000000";
		ram_buffer(5355) := X"00000000";
		ram_buffer(5356) := X"00000000";
		ram_buffer(5357) := X"00000000";
		ram_buffer(5358) := X"00000000";
		ram_buffer(5359) := X"00000000";
		ram_buffer(5360) := X"00000000";
		ram_buffer(5361) := X"00000000";
		ram_buffer(5362) := X"00000000";
		ram_buffer(5363) := X"00000000";
		ram_buffer(5364) := X"00000000";
		ram_buffer(5365) := X"00000000";
		ram_buffer(5366) := X"00000000";
		ram_buffer(5367) := X"00000000";
		ram_buffer(5368) := X"00000000";
		ram_buffer(5369) := X"00000000";
		ram_buffer(5370) := X"00000000";
		ram_buffer(5371) := X"00000000";
		ram_buffer(5372) := X"00000000";
		ram_buffer(5373) := X"00000000";
		ram_buffer(5374) := X"00000000";
		ram_buffer(5375) := X"00000000";
		ram_buffer(5376) := X"00000000";
		ram_buffer(5377) := X"00000000";
		ram_buffer(5378) := X"00000000";
		ram_buffer(5379) := X"00000000";
		ram_buffer(5380) := X"00000000";
		ram_buffer(5381) := X"00000000";
		ram_buffer(5382) := X"00000000";
		ram_buffer(5383) := X"00000000";
		ram_buffer(5384) := X"00000000";
		ram_buffer(5385) := X"00000000";
		ram_buffer(5386) := X"00000000";
		ram_buffer(5387) := X"00000000";
		ram_buffer(5388) := X"00000000";
		ram_buffer(5389) := X"00000000";
		ram_buffer(5390) := X"00000000";
		ram_buffer(5391) := X"00000000";
		ram_buffer(5392) := X"00000000";
		ram_buffer(5393) := X"00000000";
		ram_buffer(5394) := X"00000000";
		ram_buffer(5395) := X"00000000";
		ram_buffer(5396) := X"00000000";
		ram_buffer(5397) := X"00000000";
		ram_buffer(5398) := X"00000000";
		ram_buffer(5399) := X"00000000";
		ram_buffer(5400) := X"00000000";
		ram_buffer(5401) := X"00000000";
		ram_buffer(5402) := X"00000000";
		ram_buffer(5403) := X"00000000";
		ram_buffer(5404) := X"00000000";
		ram_buffer(5405) := X"00000000";
		ram_buffer(5406) := X"00000000";
		ram_buffer(5407) := X"00000000";
		ram_buffer(5408) := X"00000000";
		ram_buffer(5409) := X"00000000";
		ram_buffer(5410) := X"00000000";
		ram_buffer(5411) := X"00000000";
		ram_buffer(5412) := X"00000000";
		ram_buffer(5413) := X"00000000";
		ram_buffer(5414) := X"00000000";
		ram_buffer(5415) := X"00000000";
		ram_buffer(5416) := X"00000000";
		ram_buffer(5417) := X"00000000";
		ram_buffer(5418) := X"00000000";
		ram_buffer(5419) := X"00000000";
		ram_buffer(5420) := X"00000000";
		ram_buffer(5421) := X"00000000";
		ram_buffer(5422) := X"00000000";
		ram_buffer(5423) := X"00000000";
		ram_buffer(5424) := X"00000000";
		ram_buffer(5425) := X"00000000";
		ram_buffer(5426) := X"00000000";
		ram_buffer(5427) := X"00000000";
		ram_buffer(5428) := X"00000000";
		ram_buffer(5429) := X"00000000";
		ram_buffer(5430) := X"00000000";
		ram_buffer(5431) := X"00000000";
		ram_buffer(5432) := X"00000000";
		ram_buffer(5433) := X"00000000";
		ram_buffer(5434) := X"00000000";
		ram_buffer(5435) := X"00000000";
		ram_buffer(5436) := X"00000000";
		ram_buffer(5437) := X"00000000";
		ram_buffer(5438) := X"00000000";
		ram_buffer(5439) := X"00000000";
		ram_buffer(5440) := X"00000000";
		ram_buffer(5441) := X"00000000";
		ram_buffer(5442) := X"00000000";
		ram_buffer(5443) := X"00000000";
		ram_buffer(5444) := X"00000000";
		ram_buffer(5445) := X"00000000";
		ram_buffer(5446) := X"00000000";
		ram_buffer(5447) := X"00000000";
		ram_buffer(5448) := X"00000000";
		ram_buffer(5449) := X"00000000";
		ram_buffer(5450) := X"00000000";
		ram_buffer(5451) := X"00000000";
		ram_buffer(5452) := X"00000000";
		ram_buffer(5453) := X"00000000";
		ram_buffer(5454) := X"00000000";
		ram_buffer(5455) := X"00000000";
		ram_buffer(5456) := X"00000000";
		ram_buffer(5457) := X"00000000";
		ram_buffer(5458) := X"00000000";
		ram_buffer(5459) := X"00000000";
		ram_buffer(5460) := X"00000000";
		ram_buffer(5461) := X"00000000";
		ram_buffer(5462) := X"00000000";
		ram_buffer(5463) := X"00000000";
		ram_buffer(5464) := X"00000000";
		ram_buffer(5465) := X"00000000";
		ram_buffer(5466) := X"00000000";
		ram_buffer(5467) := X"00000000";
		ram_buffer(5468) := X"00000000";
		ram_buffer(5469) := X"00000000";
		ram_buffer(5470) := X"00000000";
		ram_buffer(5471) := X"00000000";
		ram_buffer(5472) := X"00000000";
		ram_buffer(5473) := X"00000000";
		ram_buffer(5474) := X"00000000";
		ram_buffer(5475) := X"00000000";
		ram_buffer(5476) := X"00000000";
		ram_buffer(5477) := X"00000000";
		ram_buffer(5478) := X"00000000";
		ram_buffer(5479) := X"00000000";
		ram_buffer(5480) := X"00000000";
		ram_buffer(5481) := X"00000000";
		ram_buffer(5482) := X"00000000";
		ram_buffer(5483) := X"00000000";
		ram_buffer(5484) := X"00000000";
		ram_buffer(5485) := X"00000000";
		ram_buffer(5486) := X"00000000";
		ram_buffer(5487) := X"00000000";
		ram_buffer(5488) := X"00000000";
		ram_buffer(5489) := X"00000000";
		ram_buffer(5490) := X"00000000";
		ram_buffer(5491) := X"00000000";
		ram_buffer(5492) := X"00000000";
		ram_buffer(5493) := X"00000000";
		ram_buffer(5494) := X"00000000";
		ram_buffer(5495) := X"00000000";
		ram_buffer(5496) := X"00000000";
		ram_buffer(5497) := X"00000000";
		ram_buffer(5498) := X"00000000";
		ram_buffer(5499) := X"00000000";
		ram_buffer(5500) := X"00000000";
		ram_buffer(5501) := X"00000000";
		ram_buffer(5502) := X"00000000";
		ram_buffer(5503) := X"00000000";
		ram_buffer(5504) := X"00000000";
		ram_buffer(5505) := X"00000000";
		ram_buffer(5506) := X"00000000";
		ram_buffer(5507) := X"00000000";
		ram_buffer(5508) := X"00000000";
		ram_buffer(5509) := X"00000000";
		ram_buffer(5510) := X"00000000";
		ram_buffer(5511) := X"00000000";
		ram_buffer(5512) := X"00000000";
		ram_buffer(5513) := X"00000000";
		ram_buffer(5514) := X"00000000";
		ram_buffer(5515) := X"00000000";
		ram_buffer(5516) := X"00000000";
		ram_buffer(5517) := X"00000000";
		ram_buffer(5518) := X"00000000";
		ram_buffer(5519) := X"00000000";
		ram_buffer(5520) := X"00000000";
		ram_buffer(5521) := X"00000000";
		ram_buffer(5522) := X"00000000";
		ram_buffer(5523) := X"00000000";
		ram_buffer(5524) := X"00000000";
		ram_buffer(5525) := X"00000000";
		ram_buffer(5526) := X"00000000";
		ram_buffer(5527) := X"00000000";
		ram_buffer(5528) := X"00000000";
		ram_buffer(5529) := X"00000000";
		ram_buffer(5530) := X"00000000";
		ram_buffer(5531) := X"00000000";
		ram_buffer(5532) := X"00000000";
		ram_buffer(5533) := X"00000000";
		ram_buffer(5534) := X"00000000";
		ram_buffer(5535) := X"00000000";
		ram_buffer(5536) := X"00000000";
		ram_buffer(5537) := X"00000000";
		ram_buffer(5538) := X"00000000";
		ram_buffer(5539) := X"00000000";
		ram_buffer(5540) := X"00000000";
		ram_buffer(5541) := X"00000000";
		ram_buffer(5542) := X"00000000";
		ram_buffer(5543) := X"00000000";
		ram_buffer(5544) := X"00000000";
		ram_buffer(5545) := X"00000000";
		ram_buffer(5546) := X"00000000";
		ram_buffer(5547) := X"00000000";
		ram_buffer(5548) := X"00000000";
		ram_buffer(5549) := X"00000000";
		ram_buffer(5550) := X"00000000";
		ram_buffer(5551) := X"00000000";
		ram_buffer(5552) := X"00000000";
		ram_buffer(5553) := X"00000000";
		ram_buffer(5554) := X"00000000";
		ram_buffer(5555) := X"00000000";
		ram_buffer(5556) := X"00000000";
		ram_buffer(5557) := X"00000000";
		ram_buffer(5558) := X"00000000";
		ram_buffer(5559) := X"00000000";
		ram_buffer(5560) := X"00000000";
		ram_buffer(5561) := X"00000000";
		ram_buffer(5562) := X"00000000";
		ram_buffer(5563) := X"00000000";
		ram_buffer(5564) := X"00000000";
		ram_buffer(5565) := X"00000000";
		ram_buffer(5566) := X"00000000";
		ram_buffer(5567) := X"00000000";
		ram_buffer(5568) := X"00000000";
		ram_buffer(5569) := X"00000000";
		ram_buffer(5570) := X"00000000";
		ram_buffer(5571) := X"00000000";
		ram_buffer(5572) := X"00000000";
		ram_buffer(5573) := X"00000000";
		ram_buffer(5574) := X"00000000";
		ram_buffer(5575) := X"00000000";
		ram_buffer(5576) := X"00000000";
		ram_buffer(5577) := X"00000000";
		ram_buffer(5578) := X"00000000";
		ram_buffer(5579) := X"00000000";
		ram_buffer(5580) := X"00000000";
		ram_buffer(5581) := X"00000000";
		ram_buffer(5582) := X"00000000";
		ram_buffer(5583) := X"00000000";
		ram_buffer(5584) := X"00000000";
		ram_buffer(5585) := X"00000000";
		ram_buffer(5586) := X"00000000";
		ram_buffer(5587) := X"00000000";
		ram_buffer(5588) := X"00000000";
		ram_buffer(5589) := X"00000000";
		ram_buffer(5590) := X"00000000";
		ram_buffer(5591) := X"00000000";
		ram_buffer(5592) := X"00000000";
		ram_buffer(5593) := X"00000000";
		ram_buffer(5594) := X"00000000";
		ram_buffer(5595) := X"00000000";
		ram_buffer(5596) := X"00000000";
		ram_buffer(5597) := X"00000000";
		ram_buffer(5598) := X"00000000";
		ram_buffer(5599) := X"00000000";
		ram_buffer(5600) := X"00000000";
		ram_buffer(5601) := X"00000000";
		ram_buffer(5602) := X"00000000";
		ram_buffer(5603) := X"00000000";
		ram_buffer(5604) := X"00000000";
		ram_buffer(5605) := X"00000000";
		ram_buffer(5606) := X"00000000";
		ram_buffer(5607) := X"00000000";
		ram_buffer(5608) := X"00000000";
		ram_buffer(5609) := X"00000000";
		ram_buffer(5610) := X"00000000";
		ram_buffer(5611) := X"00000000";
		ram_buffer(5612) := X"00000000";
		ram_buffer(5613) := X"00000000";
		ram_buffer(5614) := X"00000000";
		ram_buffer(5615) := X"00000000";
		ram_buffer(5616) := X"00000000";
		ram_buffer(5617) := X"00000000";
		ram_buffer(5618) := X"00000000";
		ram_buffer(5619) := X"00000000";
		ram_buffer(5620) := X"00000000";
		ram_buffer(5621) := X"00000000";
		ram_buffer(5622) := X"00000000";
		ram_buffer(5623) := X"00000000";
		ram_buffer(5624) := X"00000000";
		ram_buffer(5625) := X"00000000";
		ram_buffer(5626) := X"00000000";
		ram_buffer(5627) := X"00000000";
		ram_buffer(5628) := X"00000000";
		ram_buffer(5629) := X"00000000";
		ram_buffer(5630) := X"00000000";
		ram_buffer(5631) := X"00000000";
		ram_buffer(5632) := X"00000000";
		ram_buffer(5633) := X"00000000";
		ram_buffer(5634) := X"00000000";
		ram_buffer(5635) := X"00000000";
		ram_buffer(5636) := X"00000000";
		ram_buffer(5637) := X"00000000";
		ram_buffer(5638) := X"00000000";
		ram_buffer(5639) := X"00000000";
		ram_buffer(5640) := X"00000000";
		ram_buffer(5641) := X"00000000";
		ram_buffer(5642) := X"00000000";
		ram_buffer(5643) := X"00000000";
		ram_buffer(5644) := X"00000000";
		ram_buffer(5645) := X"00000000";
		ram_buffer(5646) := X"00000000";
		ram_buffer(5647) := X"00000000";
		ram_buffer(5648) := X"00000000";
		ram_buffer(5649) := X"00000000";
		ram_buffer(5650) := X"00000000";
		ram_buffer(5651) := X"00000000";
		ram_buffer(5652) := X"00000000";
		ram_buffer(5653) := X"00000000";
		ram_buffer(5654) := X"00000000";
		ram_buffer(5655) := X"00000000";
		ram_buffer(5656) := X"00000000";
		ram_buffer(5657) := X"00000000";
		ram_buffer(5658) := X"00000000";
		ram_buffer(5659) := X"00000000";
		ram_buffer(5660) := X"00000000";
		ram_buffer(5661) := X"00000000";
		ram_buffer(5662) := X"00000000";
		ram_buffer(5663) := X"00000000";
		ram_buffer(5664) := X"00000000";
		ram_buffer(5665) := X"00000000";
		ram_buffer(5666) := X"00000000";
		ram_buffer(5667) := X"00000000";
		ram_buffer(5668) := X"00000000";
		ram_buffer(5669) := X"00000000";
		ram_buffer(5670) := X"00000000";
		ram_buffer(5671) := X"00000000";
		ram_buffer(5672) := X"00000000";
		ram_buffer(5673) := X"00000000";
		ram_buffer(5674) := X"00000000";
		ram_buffer(5675) := X"00000000";
		ram_buffer(5676) := X"00000000";
		ram_buffer(5677) := X"00000000";
		ram_buffer(5678) := X"00000000";
		ram_buffer(5679) := X"00000000";
		ram_buffer(5680) := X"00000000";
		ram_buffer(5681) := X"00000000";
		ram_buffer(5682) := X"00000000";
		ram_buffer(5683) := X"00000000";
		ram_buffer(5684) := X"00000000";
		ram_buffer(5685) := X"00000000";
		ram_buffer(5686) := X"00000000";
		ram_buffer(5687) := X"00000000";
		ram_buffer(5688) := X"00000000";
		ram_buffer(5689) := X"00000000";
		ram_buffer(5690) := X"00000000";
		ram_buffer(5691) := X"00000000";
		ram_buffer(5692) := X"00000000";
		ram_buffer(5693) := X"00000000";
		ram_buffer(5694) := X"00000000";
		ram_buffer(5695) := X"00000000";
		ram_buffer(5696) := X"00000000";
		ram_buffer(5697) := X"00000000";
		ram_buffer(5698) := X"00000000";
		ram_buffer(5699) := X"00000000";
		ram_buffer(5700) := X"00000000";
		ram_buffer(5701) := X"00000000";
		ram_buffer(5702) := X"00000000";
		ram_buffer(5703) := X"00000000";
		ram_buffer(5704) := X"00000000";
		ram_buffer(5705) := X"00000000";
		ram_buffer(5706) := X"00000000";
		ram_buffer(5707) := X"00000000";
		ram_buffer(5708) := X"00000000";
		ram_buffer(5709) := X"00000000";
		ram_buffer(5710) := X"00000000";
		ram_buffer(5711) := X"00000000";
		ram_buffer(5712) := X"00000000";
		ram_buffer(5713) := X"00000000";
		ram_buffer(5714) := X"00000000";
		ram_buffer(5715) := X"00000000";
		ram_buffer(5716) := X"00000000";
		ram_buffer(5717) := X"00000000";
		ram_buffer(5718) := X"00000000";
		ram_buffer(5719) := X"00000000";
		ram_buffer(5720) := X"00000000";
		ram_buffer(5721) := X"00000000";
		ram_buffer(5722) := X"00000000";
		ram_buffer(5723) := X"00000000";
		ram_buffer(5724) := X"00000000";
		ram_buffer(5725) := X"00000000";
		ram_buffer(5726) := X"00000000";
		ram_buffer(5727) := X"00000000";
		ram_buffer(5728) := X"00000000";
		ram_buffer(5729) := X"00000000";
		ram_buffer(5730) := X"00000000";
		ram_buffer(5731) := X"00000000";
		ram_buffer(5732) := X"00000000";
		ram_buffer(5733) := X"00000000";
		ram_buffer(5734) := X"00000000";
		ram_buffer(5735) := X"00000000";
		ram_buffer(5736) := X"00000000";
		ram_buffer(5737) := X"00000000";
		ram_buffer(5738) := X"00000000";
		ram_buffer(5739) := X"00000000";
		ram_buffer(5740) := X"00000000";
		ram_buffer(5741) := X"00000000";
		ram_buffer(5742) := X"00000000";
		ram_buffer(5743) := X"00000000";
		ram_buffer(5744) := X"00000000";
		ram_buffer(5745) := X"00000000";
		ram_buffer(5746) := X"00000000";
		ram_buffer(5747) := X"00000000";
		ram_buffer(5748) := X"00000000";
		ram_buffer(5749) := X"00000000";
		ram_buffer(5750) := X"00000000";
		ram_buffer(5751) := X"00000000";
		ram_buffer(5752) := X"00000000";
		ram_buffer(5753) := X"00000000";
		ram_buffer(5754) := X"00000000";
		ram_buffer(5755) := X"00000000";
		ram_buffer(5756) := X"00000000";
		ram_buffer(5757) := X"00000000";
		ram_buffer(5758) := X"00000000";
		ram_buffer(5759) := X"00000000";
		ram_buffer(5760) := X"00000000";
		ram_buffer(5761) := X"00000000";
		ram_buffer(5762) := X"00000000";
		ram_buffer(5763) := X"00000000";
		ram_buffer(5764) := X"00000000";
		ram_buffer(5765) := X"00000000";
		ram_buffer(5766) := X"00000000";
		ram_buffer(5767) := X"00000000";
		ram_buffer(5768) := X"00000000";
		ram_buffer(5769) := X"00000000";
		ram_buffer(5770) := X"00000000";
		ram_buffer(5771) := X"00000000";
		ram_buffer(5772) := X"00000000";
		ram_buffer(5773) := X"00000000";
		ram_buffer(5774) := X"00000000";
		ram_buffer(5775) := X"00000000";
		ram_buffer(5776) := X"00000000";
		ram_buffer(5777) := X"00000000";
		ram_buffer(5778) := X"00000000";
		ram_buffer(5779) := X"00000000";
		ram_buffer(5780) := X"00000000";
		ram_buffer(5781) := X"00000000";
		ram_buffer(5782) := X"00000000";
		ram_buffer(5783) := X"00000000";
		ram_buffer(5784) := X"00000000";
		ram_buffer(5785) := X"00000000";
		ram_buffer(5786) := X"00000000";
		ram_buffer(5787) := X"00000000";
		ram_buffer(5788) := X"00000000";
		ram_buffer(5789) := X"00000000";
		ram_buffer(5790) := X"00000000";
		ram_buffer(5791) := X"00000000";
		ram_buffer(5792) := X"00000000";
		ram_buffer(5793) := X"00000000";
		ram_buffer(5794) := X"00000000";
		ram_buffer(5795) := X"00000000";
		ram_buffer(5796) := X"00000000";
		ram_buffer(5797) := X"00000000";
		ram_buffer(5798) := X"00000000";
		ram_buffer(5799) := X"00000000";
		ram_buffer(5800) := X"00000000";
		ram_buffer(5801) := X"00000000";
		ram_buffer(5802) := X"00000000";
		ram_buffer(5803) := X"00000000";
		ram_buffer(5804) := X"00000000";
		ram_buffer(5805) := X"00000000";
		ram_buffer(5806) := X"00000000";
		ram_buffer(5807) := X"00000000";
		ram_buffer(5808) := X"00000000";
		ram_buffer(5809) := X"00000000";
		ram_buffer(5810) := X"00000000";
		ram_buffer(5811) := X"00000000";
		ram_buffer(5812) := X"00000000";
		ram_buffer(5813) := X"00000000";
		ram_buffer(5814) := X"00000000";
		ram_buffer(5815) := X"00000000";
		ram_buffer(5816) := X"00000000";
		ram_buffer(5817) := X"00000000";
		ram_buffer(5818) := X"00000000";
		ram_buffer(5819) := X"00000000";
		ram_buffer(5820) := X"00000000";
		ram_buffer(5821) := X"00000000";
		ram_buffer(5822) := X"00000000";
		ram_buffer(5823) := X"00000000";
		ram_buffer(5824) := X"00000000";
		ram_buffer(5825) := X"00000000";
		ram_buffer(5826) := X"00000000";
		ram_buffer(5827) := X"00000000";
		ram_buffer(5828) := X"00000000";
		ram_buffer(5829) := X"00000000";
		ram_buffer(5830) := X"00000000";
		ram_buffer(5831) := X"00000000";
		ram_buffer(5832) := X"00000000";
		ram_buffer(5833) := X"00000000";
		ram_buffer(5834) := X"00000000";
		ram_buffer(5835) := X"00000000";
		ram_buffer(5836) := X"00000000";
		ram_buffer(5837) := X"00000000";
		ram_buffer(5838) := X"00000000";
		ram_buffer(5839) := X"00000000";
		ram_buffer(5840) := X"00000000";
		ram_buffer(5841) := X"00000000";
		ram_buffer(5842) := X"00000000";
		ram_buffer(5843) := X"00000000";
		ram_buffer(5844) := X"00000000";
		ram_buffer(5845) := X"00000000";
		ram_buffer(5846) := X"00000000";
		ram_buffer(5847) := X"00000000";
		ram_buffer(5848) := X"00000000";
		ram_buffer(5849) := X"00000000";
		ram_buffer(5850) := X"00000000";
		ram_buffer(5851) := X"00000000";
		ram_buffer(5852) := X"00000000";
		ram_buffer(5853) := X"00000000";
		ram_buffer(5854) := X"00000000";
		ram_buffer(5855) := X"00000000";
		ram_buffer(5856) := X"00000000";
		ram_buffer(5857) := X"00000000";
		ram_buffer(5858) := X"00000000";
		ram_buffer(5859) := X"00000000";
		ram_buffer(5860) := X"00000000";
		ram_buffer(5861) := X"00000000";
		ram_buffer(5862) := X"00000000";
		ram_buffer(5863) := X"00000000";
		ram_buffer(5864) := X"00000000";
		ram_buffer(5865) := X"00000000";
		ram_buffer(5866) := X"00000000";
		ram_buffer(5867) := X"00000000";
		ram_buffer(5868) := X"00000000";
		ram_buffer(5869) := X"00000000";
		ram_buffer(5870) := X"00000000";
		ram_buffer(5871) := X"00000000";
		ram_buffer(5872) := X"00000000";
		ram_buffer(5873) := X"00000000";
		ram_buffer(5874) := X"00000000";
		ram_buffer(5875) := X"00000000";
		ram_buffer(5876) := X"00000000";
		ram_buffer(5877) := X"00000000";
		ram_buffer(5878) := X"00000000";
		ram_buffer(5879) := X"00000000";
		ram_buffer(5880) := X"00000000";
		ram_buffer(5881) := X"00000000";
		ram_buffer(5882) := X"00000000";
		ram_buffer(5883) := X"00000000";
		ram_buffer(5884) := X"00000000";
		ram_buffer(5885) := X"00000000";
		ram_buffer(5886) := X"00000000";
		ram_buffer(5887) := X"00000000";
		ram_buffer(5888) := X"00000000";
		ram_buffer(5889) := X"00000000";
		ram_buffer(5890) := X"00000000";
		ram_buffer(5891) := X"00000000";
		ram_buffer(5892) := X"00000000";
		ram_buffer(5893) := X"00000000";
		ram_buffer(5894) := X"00000000";
		ram_buffer(5895) := X"00000000";
		ram_buffer(5896) := X"00000000";
		ram_buffer(5897) := X"00000000";
		ram_buffer(5898) := X"00000000";
		ram_buffer(5899) := X"00000000";
		ram_buffer(5900) := X"00000000";
		ram_buffer(5901) := X"00000000";
		ram_buffer(5902) := X"00000000";
		ram_buffer(5903) := X"00000000";
		ram_buffer(5904) := X"00000000";
		ram_buffer(5905) := X"00000000";
		ram_buffer(5906) := X"00000000";
		ram_buffer(5907) := X"00000000";
		ram_buffer(5908) := X"00000000";
		ram_buffer(5909) := X"00000000";
		ram_buffer(5910) := X"00000000";
		ram_buffer(5911) := X"00000000";
		ram_buffer(5912) := X"00000000";
		ram_buffer(5913) := X"00000000";
		ram_buffer(5914) := X"00000000";
		ram_buffer(5915) := X"00000000";
		ram_buffer(5916) := X"00000000";
		ram_buffer(5917) := X"00000000";
		ram_buffer(5918) := X"00000000";
		ram_buffer(5919) := X"00000000";
		ram_buffer(5920) := X"00000000";
		ram_buffer(5921) := X"00000000";
		ram_buffer(5922) := X"00000000";
		ram_buffer(5923) := X"00000000";
		ram_buffer(5924) := X"00000000";
		ram_buffer(5925) := X"00000000";
		ram_buffer(5926) := X"00000000";
		ram_buffer(5927) := X"00000000";
		ram_buffer(5928) := X"00000000";
		ram_buffer(5929) := X"00000000";
		ram_buffer(5930) := X"00000000";
		ram_buffer(5931) := X"00000000";
		ram_buffer(5932) := X"00000000";
		ram_buffer(5933) := X"00000000";
		ram_buffer(5934) := X"00000000";
		ram_buffer(5935) := X"00000000";
		ram_buffer(5936) := X"00000000";
		ram_buffer(5937) := X"00000000";
		ram_buffer(5938) := X"00000000";
		ram_buffer(5939) := X"00000000";
		ram_buffer(5940) := X"00000000";
		ram_buffer(5941) := X"00000000";
		ram_buffer(5942) := X"00000000";
		ram_buffer(5943) := X"00000000";
		ram_buffer(5944) := X"00000000";
		ram_buffer(5945) := X"00000000";
		ram_buffer(5946) := X"00000000";
		ram_buffer(5947) := X"00000000";
		ram_buffer(5948) := X"00000000";
		ram_buffer(5949) := X"00000000";
		ram_buffer(5950) := X"00000000";
		ram_buffer(5951) := X"00000000";
		ram_buffer(5952) := X"00000000";
		ram_buffer(5953) := X"00000000";
		ram_buffer(5954) := X"00000000";
		ram_buffer(5955) := X"00000000";
		ram_buffer(5956) := X"00000000";
		ram_buffer(5957) := X"00000000";
		ram_buffer(5958) := X"00000000";
		ram_buffer(5959) := X"00000000";
		ram_buffer(5960) := X"00000000";
		ram_buffer(5961) := X"00000000";
		ram_buffer(5962) := X"00000000";
		ram_buffer(5963) := X"00000000";
		ram_buffer(5964) := X"00000000";
		ram_buffer(5965) := X"00000000";
		ram_buffer(5966) := X"00000000";
		ram_buffer(5967) := X"00000000";
		ram_buffer(5968) := X"00000000";
		ram_buffer(5969) := X"00000000";
		ram_buffer(5970) := X"00000000";
		ram_buffer(5971) := X"00000000";
		ram_buffer(5972) := X"00000000";
		ram_buffer(5973) := X"00000000";
		ram_buffer(5974) := X"00000000";
		ram_buffer(5975) := X"00000000";
		ram_buffer(5976) := X"00000000";
		ram_buffer(5977) := X"00000000";
		ram_buffer(5978) := X"00000000";
		ram_buffer(5979) := X"00000000";
		ram_buffer(5980) := X"00000000";
		ram_buffer(5981) := X"00000000";
		ram_buffer(5982) := X"00000000";
		ram_buffer(5983) := X"00000000";
		ram_buffer(5984) := X"00000000";
		ram_buffer(5985) := X"00000000";
		ram_buffer(5986) := X"00000000";
		ram_buffer(5987) := X"00000000";
		ram_buffer(5988) := X"00000000";
		ram_buffer(5989) := X"00000000";
		ram_buffer(5990) := X"00000000";
		ram_buffer(5991) := X"00000000";
		ram_buffer(5992) := X"00000000";
		ram_buffer(5993) := X"00000000";
		ram_buffer(5994) := X"00000000";
		ram_buffer(5995) := X"00000000";
		ram_buffer(5996) := X"00000000";
		ram_buffer(5997) := X"00000000";
		ram_buffer(5998) := X"00000000";
		ram_buffer(5999) := X"00000000";
		ram_buffer(6000) := X"00000000";
		ram_buffer(6001) := X"00000000";
		ram_buffer(6002) := X"00000000";
		ram_buffer(6003) := X"00000000";
		ram_buffer(6004) := X"00000000";
		ram_buffer(6005) := X"00000000";
		ram_buffer(6006) := X"00000000";
		ram_buffer(6007) := X"00000000";
		ram_buffer(6008) := X"00000000";
		ram_buffer(6009) := X"00000000";
		ram_buffer(6010) := X"00000000";
		ram_buffer(6011) := X"00000000";
		ram_buffer(6012) := X"00000000";
		ram_buffer(6013) := X"00000000";
		ram_buffer(6014) := X"00000000";
		ram_buffer(6015) := X"00000000";
		ram_buffer(6016) := X"00000000";
		ram_buffer(6017) := X"00000000";
		ram_buffer(6018) := X"00000000";
		ram_buffer(6019) := X"00000000";
		ram_buffer(6020) := X"00000000";
		ram_buffer(6021) := X"00000000";
		ram_buffer(6022) := X"00000000";
		ram_buffer(6023) := X"00000000";
		ram_buffer(6024) := X"00000000";
		ram_buffer(6025) := X"00000000";
		ram_buffer(6026) := X"00000000";
		ram_buffer(6027) := X"00000000";
		ram_buffer(6028) := X"00000000";
		ram_buffer(6029) := X"00000000";
		ram_buffer(6030) := X"00000000";
		ram_buffer(6031) := X"00000000";
		ram_buffer(6032) := X"00000000";
		ram_buffer(6033) := X"00000000";
		ram_buffer(6034) := X"00000000";
		ram_buffer(6035) := X"00000000";
		ram_buffer(6036) := X"00000000";
		ram_buffer(6037) := X"00000000";
		ram_buffer(6038) := X"00000000";
		ram_buffer(6039) := X"00000000";
		ram_buffer(6040) := X"00000000";
		ram_buffer(6041) := X"00000000";
		ram_buffer(6042) := X"00000000";
		ram_buffer(6043) := X"00000000";
		ram_buffer(6044) := X"00000000";
		ram_buffer(6045) := X"00000000";
		ram_buffer(6046) := X"00000000";
		ram_buffer(6047) := X"00000000";
		ram_buffer(6048) := X"00000000";
		ram_buffer(6049) := X"00000000";
		ram_buffer(6050) := X"00000000";
		ram_buffer(6051) := X"00000000";
		ram_buffer(6052) := X"00000000";
		ram_buffer(6053) := X"00000000";
		ram_buffer(6054) := X"00000000";
		ram_buffer(6055) := X"00000000";
		ram_buffer(6056) := X"00000000";
		ram_buffer(6057) := X"00000000";
		ram_buffer(6058) := X"00000000";
		ram_buffer(6059) := X"00000000";
		ram_buffer(6060) := X"00000000";
		ram_buffer(6061) := X"00000000";
		ram_buffer(6062) := X"00000000";
		ram_buffer(6063) := X"00000000";
		ram_buffer(6064) := X"00000000";
		ram_buffer(6065) := X"00000000";
		ram_buffer(6066) := X"00000000";
		ram_buffer(6067) := X"00000000";
		ram_buffer(6068) := X"00000000";
		ram_buffer(6069) := X"00000000";
		ram_buffer(6070) := X"00000000";
		ram_buffer(6071) := X"00000000";
		ram_buffer(6072) := X"00000000";
		ram_buffer(6073) := X"00000000";
		ram_buffer(6074) := X"00000000";
		ram_buffer(6075) := X"00000000";
		ram_buffer(6076) := X"00000000";
		ram_buffer(6077) := X"00000000";
		ram_buffer(6078) := X"00000000";
		ram_buffer(6079) := X"00000000";
		ram_buffer(6080) := X"00000000";
		ram_buffer(6081) := X"00000000";
		ram_buffer(6082) := X"00000000";
		ram_buffer(6083) := X"00000000";
		ram_buffer(6084) := X"00000000";
		ram_buffer(6085) := X"00000000";
		ram_buffer(6086) := X"00000000";
		ram_buffer(6087) := X"00000000";
		ram_buffer(6088) := X"00000000";
		ram_buffer(6089) := X"00000000";
		ram_buffer(6090) := X"00000000";
		ram_buffer(6091) := X"00000000";
		ram_buffer(6092) := X"00000000";
		ram_buffer(6093) := X"00000000";
		ram_buffer(6094) := X"00000000";
		ram_buffer(6095) := X"00000000";
		ram_buffer(6096) := X"00000000";
		ram_buffer(6097) := X"00000000";
		ram_buffer(6098) := X"00000000";
		ram_buffer(6099) := X"00000000";
		ram_buffer(6100) := X"00000000";
		ram_buffer(6101) := X"00000000";
		ram_buffer(6102) := X"00000000";
		ram_buffer(6103) := X"00000000";
		ram_buffer(6104) := X"00000000";
		ram_buffer(6105) := X"00000000";
		ram_buffer(6106) := X"00000000";
		ram_buffer(6107) := X"00000000";
		ram_buffer(6108) := X"00000000";
		ram_buffer(6109) := X"00000000";
		ram_buffer(6110) := X"00000000";
		ram_buffer(6111) := X"00000000";
		ram_buffer(6112) := X"00000000";
		ram_buffer(6113) := X"00000000";
		ram_buffer(6114) := X"00000000";
		ram_buffer(6115) := X"00000000";
		ram_buffer(6116) := X"00000000";
		ram_buffer(6117) := X"00000000";
		ram_buffer(6118) := X"00000000";
		ram_buffer(6119) := X"00000000";
		ram_buffer(6120) := X"00000000";
		ram_buffer(6121) := X"00000000";
		ram_buffer(6122) := X"00000000";
		ram_buffer(6123) := X"00000000";
		ram_buffer(6124) := X"00000000";
		ram_buffer(6125) := X"00000000";
		ram_buffer(6126) := X"00000000";
		ram_buffer(6127) := X"00000000";
		ram_buffer(6128) := X"00000000";
		ram_buffer(6129) := X"00000000";
		ram_buffer(6130) := X"00000000";
		ram_buffer(6131) := X"00000000";
		ram_buffer(6132) := X"00000000";
		ram_buffer(6133) := X"00000000";
		ram_buffer(6134) := X"00000000";
		ram_buffer(6135) := X"00000000";
		ram_buffer(6136) := X"00000000";
		ram_buffer(6137) := X"00000000";
		ram_buffer(6138) := X"00000000";
		ram_buffer(6139) := X"00000000";
		ram_buffer(6140) := X"00000000";
		ram_buffer(6141) := X"00000000";
		ram_buffer(6142) := X"00000000";
		ram_buffer(6143) := X"00000000";
		ram_buffer(6144) := X"00000000";
		ram_buffer(6145) := X"00000000";
		ram_buffer(6146) := X"00000000";
		ram_buffer(6147) := X"00000000";
		ram_buffer(6148) := X"00000000";
		ram_buffer(6149) := X"00000000";
		ram_buffer(6150) := X"00000000";
		ram_buffer(6151) := X"00000000";
		ram_buffer(6152) := X"00000000";
		ram_buffer(6153) := X"00000000";
		ram_buffer(6154) := X"00000000";
		ram_buffer(6155) := X"00000000";
		ram_buffer(6156) := X"00000000";
		ram_buffer(6157) := X"00000000";
		ram_buffer(6158) := X"00000000";
		ram_buffer(6159) := X"00000000";
		ram_buffer(6160) := X"00000000";
		ram_buffer(6161) := X"00000000";
		ram_buffer(6162) := X"00000000";
		ram_buffer(6163) := X"00000000";
		ram_buffer(6164) := X"00000000";
		ram_buffer(6165) := X"00000000";
		ram_buffer(6166) := X"00000000";
		ram_buffer(6167) := X"00000000";
		ram_buffer(6168) := X"00000000";
		ram_buffer(6169) := X"00000000";
		ram_buffer(6170) := X"00000000";
		ram_buffer(6171) := X"00000000";
		ram_buffer(6172) := X"00000000";
		ram_buffer(6173) := X"00000000";
		ram_buffer(6174) := X"00000000";
		ram_buffer(6175) := X"00000000";
		ram_buffer(6176) := X"00000000";
		ram_buffer(6177) := X"00000000";
		ram_buffer(6178) := X"00000000";
		ram_buffer(6179) := X"00000000";
		ram_buffer(6180) := X"00000000";
		ram_buffer(6181) := X"00000000";
		ram_buffer(6182) := X"00000000";
		ram_buffer(6183) := X"00000000";
		ram_buffer(6184) := X"00000000";
		ram_buffer(6185) := X"00000000";
		ram_buffer(6186) := X"00000000";
		ram_buffer(6187) := X"00000000";
		ram_buffer(6188) := X"00000000";
		ram_buffer(6189) := X"00000000";
		ram_buffer(6190) := X"00000000";
		ram_buffer(6191) := X"00000000";
		ram_buffer(6192) := X"00000000";
		ram_buffer(6193) := X"00000000";
		ram_buffer(6194) := X"00000000";
		ram_buffer(6195) := X"00000000";
		ram_buffer(6196) := X"00000000";
		ram_buffer(6197) := X"00000000";
		ram_buffer(6198) := X"00000000";
		ram_buffer(6199) := X"00000000";
		ram_buffer(6200) := X"00000000";
		ram_buffer(6201) := X"00000000";
		ram_buffer(6202) := X"00000000";
		ram_buffer(6203) := X"00000000";
		ram_buffer(6204) := X"00000000";
		ram_buffer(6205) := X"00000000";
		ram_buffer(6206) := X"00000000";
		ram_buffer(6207) := X"00000000";
		ram_buffer(6208) := X"00000000";
		ram_buffer(6209) := X"00000000";
		ram_buffer(6210) := X"00000000";
		ram_buffer(6211) := X"00000000";
		ram_buffer(6212) := X"00000000";
		ram_buffer(6213) := X"00000000";
		ram_buffer(6214) := X"00000000";
		ram_buffer(6215) := X"00000000";
		ram_buffer(6216) := X"00000000";
		ram_buffer(6217) := X"00000000";
		ram_buffer(6218) := X"00000000";
		ram_buffer(6219) := X"00000000";
		ram_buffer(6220) := X"00000000";
		ram_buffer(6221) := X"00000000";
		ram_buffer(6222) := X"00000000";
		ram_buffer(6223) := X"00000000";
		ram_buffer(6224) := X"00000000";
		ram_buffer(6225) := X"00000000";
		ram_buffer(6226) := X"00000000";
		ram_buffer(6227) := X"00000000";
		ram_buffer(6228) := X"00000000";
		ram_buffer(6229) := X"00000000";
		ram_buffer(6230) := X"00000000";
		ram_buffer(6231) := X"00000000";
		ram_buffer(6232) := X"00000000";
		ram_buffer(6233) := X"00000000";
		ram_buffer(6234) := X"00000000";
		ram_buffer(6235) := X"00000000";
		ram_buffer(6236) := X"00000000";
		ram_buffer(6237) := X"00000000";
		ram_buffer(6238) := X"00000000";
		ram_buffer(6239) := X"00000000";
		ram_buffer(6240) := X"00000000";
		ram_buffer(6241) := X"00000000";
		ram_buffer(6242) := X"00000000";
		ram_buffer(6243) := X"00000000";
		ram_buffer(6244) := X"00000000";
		ram_buffer(6245) := X"00000000";
		ram_buffer(6246) := X"00000000";
		ram_buffer(6247) := X"00000000";
		ram_buffer(6248) := X"00000000";
		ram_buffer(6249) := X"00000000";
		ram_buffer(6250) := X"00000000";
		ram_buffer(6251) := X"00000000";
		ram_buffer(6252) := X"00000000";
		ram_buffer(6253) := X"00000000";
		ram_buffer(6254) := X"00000000";
		ram_buffer(6255) := X"00000000";
		ram_buffer(6256) := X"00000000";
		ram_buffer(6257) := X"00000000";
		ram_buffer(6258) := X"00000000";
		ram_buffer(6259) := X"00000000";
		ram_buffer(6260) := X"00000000";
		ram_buffer(6261) := X"00000000";
		ram_buffer(6262) := X"00000000";
		ram_buffer(6263) := X"00000000";
		ram_buffer(6264) := X"00000000";
		ram_buffer(6265) := X"00000000";
		ram_buffer(6266) := X"00000000";
		ram_buffer(6267) := X"00000000";
		ram_buffer(6268) := X"00000000";
		ram_buffer(6269) := X"00000000";
		ram_buffer(6270) := X"00000000";
		ram_buffer(6271) := X"00000000";
		ram_buffer(6272) := X"00000000";
		ram_buffer(6273) := X"00000000";
		ram_buffer(6274) := X"00000000";
		ram_buffer(6275) := X"00000000";
		ram_buffer(6276) := X"00000000";
		ram_buffer(6277) := X"00000000";
		ram_buffer(6278) := X"00000000";
		ram_buffer(6279) := X"00000000";
		ram_buffer(6280) := X"00000000";
		ram_buffer(6281) := X"00000000";
		ram_buffer(6282) := X"00000000";
		ram_buffer(6283) := X"00000000";
		ram_buffer(6284) := X"00000000";
		ram_buffer(6285) := X"00000000";
		ram_buffer(6286) := X"00000000";
		ram_buffer(6287) := X"00000000";
		ram_buffer(6288) := X"00000000";
		ram_buffer(6289) := X"00000000";
		ram_buffer(6290) := X"00000000";
		ram_buffer(6291) := X"00000000";
		ram_buffer(6292) := X"00000000";
		ram_buffer(6293) := X"00000000";
		ram_buffer(6294) := X"00000000";
		ram_buffer(6295) := X"00000000";
		ram_buffer(6296) := X"00000000";
		ram_buffer(6297) := X"00000000";
		ram_buffer(6298) := X"00000000";
		ram_buffer(6299) := X"00000000";
		ram_buffer(6300) := X"00000000";
		ram_buffer(6301) := X"00000000";
		ram_buffer(6302) := X"00000000";
		ram_buffer(6303) := X"00000000";
		ram_buffer(6304) := X"00000000";
		ram_buffer(6305) := X"00000000";
		ram_buffer(6306) := X"00000000";
		ram_buffer(6307) := X"00000000";
		ram_buffer(6308) := X"00000000";
		ram_buffer(6309) := X"00000000";
		ram_buffer(6310) := X"00000000";
		ram_buffer(6311) := X"00000000";
		ram_buffer(6312) := X"00000000";
		ram_buffer(6313) := X"00000000";
		ram_buffer(6314) := X"00000000";
		ram_buffer(6315) := X"00000000";
		ram_buffer(6316) := X"00000000";
		ram_buffer(6317) := X"00000000";
		ram_buffer(6318) := X"00000000";
		ram_buffer(6319) := X"00000000";
		ram_buffer(6320) := X"00000000";
		ram_buffer(6321) := X"00000000";
		ram_buffer(6322) := X"00000000";
		ram_buffer(6323) := X"00000000";
		ram_buffer(6324) := X"00000000";
		ram_buffer(6325) := X"00000000";
		ram_buffer(6326) := X"00000000";
		ram_buffer(6327) := X"00000000";
		ram_buffer(6328) := X"00000000";
		ram_buffer(6329) := X"00000000";
		ram_buffer(6330) := X"00000000";
		ram_buffer(6331) := X"00000000";
		ram_buffer(6332) := X"00000000";
		ram_buffer(6333) := X"00000000";
		ram_buffer(6334) := X"00000000";
		ram_buffer(6335) := X"00000000";
		ram_buffer(6336) := X"00000000";
		ram_buffer(6337) := X"00000000";
		ram_buffer(6338) := X"00000000";
		ram_buffer(6339) := X"00000000";
		ram_buffer(6340) := X"00000000";
		ram_buffer(6341) := X"00000000";
		ram_buffer(6342) := X"00000000";
		ram_buffer(6343) := X"00000000";
		ram_buffer(6344) := X"00000000";
		ram_buffer(6345) := X"00000000";
		ram_buffer(6346) := X"00000000";
		ram_buffer(6347) := X"00000000";
		ram_buffer(6348) := X"00000000";
		ram_buffer(6349) := X"00000000";
		ram_buffer(6350) := X"00000000";
		ram_buffer(6351) := X"00000000";
		ram_buffer(6352) := X"00000000";
		ram_buffer(6353) := X"00000000";
		ram_buffer(6354) := X"00000000";
		ram_buffer(6355) := X"00000000";
		ram_buffer(6356) := X"00000000";
		ram_buffer(6357) := X"00000000";
		ram_buffer(6358) := X"00000000";
		ram_buffer(6359) := X"00000000";
		ram_buffer(6360) := X"00000000";
		ram_buffer(6361) := X"00000000";
		ram_buffer(6362) := X"00000000";
		ram_buffer(6363) := X"00000000";
		ram_buffer(6364) := X"00000000";
		ram_buffer(6365) := X"00000000";
		ram_buffer(6366) := X"00000000";
		ram_buffer(6367) := X"00000000";
		ram_buffer(6368) := X"00000000";
		ram_buffer(6369) := X"00000000";
		ram_buffer(6370) := X"00000000";
		ram_buffer(6371) := X"00000000";
		ram_buffer(6372) := X"00000000";
		ram_buffer(6373) := X"00000000";
		ram_buffer(6374) := X"00000000";
		ram_buffer(6375) := X"00000000";
		ram_buffer(6376) := X"00000000";
		ram_buffer(6377) := X"00000000";
		ram_buffer(6378) := X"00000000";
		ram_buffer(6379) := X"00000000";
		ram_buffer(6380) := X"00000000";
		ram_buffer(6381) := X"00000000";
		ram_buffer(6382) := X"00000000";
		ram_buffer(6383) := X"00000000";
		ram_buffer(6384) := X"00000000";
		ram_buffer(6385) := X"00000000";
		ram_buffer(6386) := X"00000000";
		ram_buffer(6387) := X"00000000";
		ram_buffer(6388) := X"00000000";
		ram_buffer(6389) := X"00000000";
		ram_buffer(6390) := X"00000000";
		ram_buffer(6391) := X"00000000";
		ram_buffer(6392) := X"00000000";
		ram_buffer(6393) := X"00000000";
		ram_buffer(6394) := X"00000000";
		ram_buffer(6395) := X"00000000";
		ram_buffer(6396) := X"00000000";
		ram_buffer(6397) := X"00000000";
		ram_buffer(6398) := X"00000000";
		ram_buffer(6399) := X"00000000";
		ram_buffer(6400) := X"00000000";
		ram_buffer(6401) := X"00000000";
		ram_buffer(6402) := X"00000000";
		ram_buffer(6403) := X"00000000";
		ram_buffer(6404) := X"00000000";
		ram_buffer(6405) := X"00000000";
		ram_buffer(6406) := X"00000000";
		ram_buffer(6407) := X"00000000";
		ram_buffer(6408) := X"00000000";
		ram_buffer(6409) := X"00000000";
		ram_buffer(6410) := X"00000000";
		ram_buffer(6411) := X"00000000";
		ram_buffer(6412) := X"00000000";
		ram_buffer(6413) := X"00000000";
		ram_buffer(6414) := X"00000000";
		ram_buffer(6415) := X"00000000";
		ram_buffer(6416) := X"00000000";
		ram_buffer(6417) := X"00000000";
		ram_buffer(6418) := X"00000000";
		ram_buffer(6419) := X"00000000";
		ram_buffer(6420) := X"00000000";
		ram_buffer(6421) := X"00000000";
		ram_buffer(6422) := X"00000000";
		ram_buffer(6423) := X"00000000";
		ram_buffer(6424) := X"00000000";
		ram_buffer(6425) := X"00000000";
		ram_buffer(6426) := X"00000000";
		ram_buffer(6427) := X"00000000";
		ram_buffer(6428) := X"00000000";
		ram_buffer(6429) := X"00000000";
		ram_buffer(6430) := X"00000000";
		ram_buffer(6431) := X"00000000";
		ram_buffer(6432) := X"00000000";
		ram_buffer(6433) := X"00000000";
		ram_buffer(6434) := X"00000000";
		ram_buffer(6435) := X"00000000";
		ram_buffer(6436) := X"00000000";
		ram_buffer(6437) := X"00000000";
		ram_buffer(6438) := X"00000000";
		ram_buffer(6439) := X"00000000";
		ram_buffer(6440) := X"00000000";
		ram_buffer(6441) := X"00000000";
		ram_buffer(6442) := X"00000000";
		ram_buffer(6443) := X"00000000";
		ram_buffer(6444) := X"00000000";
		ram_buffer(6445) := X"00000000";
		ram_buffer(6446) := X"00000000";
		ram_buffer(6447) := X"00000000";
		ram_buffer(6448) := X"00000000";
		ram_buffer(6449) := X"00000000";
		ram_buffer(6450) := X"00000000";
		ram_buffer(6451) := X"00000000";
		ram_buffer(6452) := X"00000000";
		ram_buffer(6453) := X"00000000";
		ram_buffer(6454) := X"00000000";
		ram_buffer(6455) := X"00000000";
		ram_buffer(6456) := X"00000000";
		ram_buffer(6457) := X"00000000";
		ram_buffer(6458) := X"00000000";
		ram_buffer(6459) := X"00000000";
		ram_buffer(6460) := X"00000000";
		ram_buffer(6461) := X"00000000";
		ram_buffer(6462) := X"00000000";
		ram_buffer(6463) := X"00000000";
		ram_buffer(6464) := X"00000000";
		ram_buffer(6465) := X"00000000";
		ram_buffer(6466) := X"00000000";
		ram_buffer(6467) := X"00000000";
		ram_buffer(6468) := X"00000000";
		ram_buffer(6469) := X"00000000";
		ram_buffer(6470) := X"00000000";
		ram_buffer(6471) := X"00000000";
		ram_buffer(6472) := X"00000000";
		ram_buffer(6473) := X"00000000";
		ram_buffer(6474) := X"00000000";
		ram_buffer(6475) := X"00000000";
		ram_buffer(6476) := X"00000000";
		ram_buffer(6477) := X"00000000";
		ram_buffer(6478) := X"00000000";
		ram_buffer(6479) := X"00000000";
		ram_buffer(6480) := X"00000000";
		ram_buffer(6481) := X"00000000";
		ram_buffer(6482) := X"00000000";
		ram_buffer(6483) := X"00000000";
		ram_buffer(6484) := X"00000000";
		ram_buffer(6485) := X"00000000";
		ram_buffer(6486) := X"00000000";
		ram_buffer(6487) := X"00000000";
		ram_buffer(6488) := X"00000000";
		ram_buffer(6489) := X"00000000";
		ram_buffer(6490) := X"00000000";
		ram_buffer(6491) := X"00000000";
		ram_buffer(6492) := X"00000000";
		ram_buffer(6493) := X"00000000";
		ram_buffer(6494) := X"00000000";
		ram_buffer(6495) := X"00000000";
		ram_buffer(6496) := X"00000000";
		ram_buffer(6497) := X"00000000";
		ram_buffer(6498) := X"00000000";
		ram_buffer(6499) := X"00000000";
		ram_buffer(6500) := X"00000000";
		ram_buffer(6501) := X"00000000";
		ram_buffer(6502) := X"00000000";
		ram_buffer(6503) := X"00000000";
		ram_buffer(6504) := X"00000000";
		ram_buffer(6505) := X"00000000";
		ram_buffer(6506) := X"00000000";
		ram_buffer(6507) := X"00000000";
		ram_buffer(6508) := X"00000000";
		ram_buffer(6509) := X"00000000";
		ram_buffer(6510) := X"00000000";
		ram_buffer(6511) := X"00000000";
		ram_buffer(6512) := X"00000000";
		ram_buffer(6513) := X"00000000";
		ram_buffer(6514) := X"00000000";
		ram_buffer(6515) := X"00000000";
		ram_buffer(6516) := X"00000000";
		ram_buffer(6517) := X"00000000";
		ram_buffer(6518) := X"00000000";
		ram_buffer(6519) := X"00000000";
		ram_buffer(6520) := X"00000000";
		ram_buffer(6521) := X"00000000";
		ram_buffer(6522) := X"00000000";
		ram_buffer(6523) := X"00000000";
		ram_buffer(6524) := X"00000000";
		ram_buffer(6525) := X"00000000";
		ram_buffer(6526) := X"00000000";
		ram_buffer(6527) := X"00000000";
		ram_buffer(6528) := X"00000000";
		ram_buffer(6529) := X"00000000";
		ram_buffer(6530) := X"00000000";
		ram_buffer(6531) := X"00000000";
		ram_buffer(6532) := X"00000000";
		ram_buffer(6533) := X"00000000";
		ram_buffer(6534) := X"00000000";
		ram_buffer(6535) := X"00000000";
		ram_buffer(6536) := X"00000000";
		ram_buffer(6537) := X"00000000";
		ram_buffer(6538) := X"00000000";
		ram_buffer(6539) := X"00000000";
		ram_buffer(6540) := X"00000000";
		ram_buffer(6541) := X"00000000";
		ram_buffer(6542) := X"00000000";
		ram_buffer(6543) := X"00000000";
		ram_buffer(6544) := X"00000000";
		ram_buffer(6545) := X"00000000";
		ram_buffer(6546) := X"00000000";
		ram_buffer(6547) := X"00000000";
		ram_buffer(6548) := X"00000000";
		ram_buffer(6549) := X"00000000";
		ram_buffer(6550) := X"00000000";
		ram_buffer(6551) := X"00000000";
		ram_buffer(6552) := X"00000000";
		ram_buffer(6553) := X"00000000";
		ram_buffer(6554) := X"00000000";
		ram_buffer(6555) := X"00000000";
		ram_buffer(6556) := X"00000000";
		ram_buffer(6557) := X"00000000";
		ram_buffer(6558) := X"00000000";
		ram_buffer(6559) := X"00000000";
		ram_buffer(6560) := X"00000000";
		ram_buffer(6561) := X"00000000";
		ram_buffer(6562) := X"00000000";
		ram_buffer(6563) := X"00000000";
		ram_buffer(6564) := X"00000000";
		ram_buffer(6565) := X"00000000";
		ram_buffer(6566) := X"00000000";
		ram_buffer(6567) := X"00000000";
		ram_buffer(6568) := X"00000000";
		ram_buffer(6569) := X"00000000";
		ram_buffer(6570) := X"00000000";
		ram_buffer(6571) := X"00000000";
		ram_buffer(6572) := X"00000000";
		ram_buffer(6573) := X"00000000";
		ram_buffer(6574) := X"00000000";
		ram_buffer(6575) := X"00000000";
		ram_buffer(6576) := X"00000000";
		ram_buffer(6577) := X"00000000";
		ram_buffer(6578) := X"00000000";
		ram_buffer(6579) := X"00000000";
		ram_buffer(6580) := X"00000000";
		ram_buffer(6581) := X"00000000";
		ram_buffer(6582) := X"00000000";
		ram_buffer(6583) := X"00000000";
		ram_buffer(6584) := X"00000000";
		ram_buffer(6585) := X"00000000";
		ram_buffer(6586) := X"00000000";
		ram_buffer(6587) := X"00000000";
		ram_buffer(6588) := X"00000000";
		ram_buffer(6589) := X"00000000";
		ram_buffer(6590) := X"00000000";
		ram_buffer(6591) := X"00000000";
		ram_buffer(6592) := X"00000000";
		ram_buffer(6593) := X"00000000";
		ram_buffer(6594) := X"00000000";
		ram_buffer(6595) := X"00000000";
		ram_buffer(6596) := X"00000000";
		ram_buffer(6597) := X"00000000";
		ram_buffer(6598) := X"00000000";
		ram_buffer(6599) := X"00000000";
		ram_buffer(6600) := X"00000000";
		ram_buffer(6601) := X"00000000";
		ram_buffer(6602) := X"00000000";
		ram_buffer(6603) := X"00000000";
		ram_buffer(6604) := X"00000000";
		ram_buffer(6605) := X"00000000";
		ram_buffer(6606) := X"00000000";
		ram_buffer(6607) := X"00000000";
		ram_buffer(6608) := X"00000000";
		ram_buffer(6609) := X"00000000";
		ram_buffer(6610) := X"00000000";
		ram_buffer(6611) := X"00000000";
		ram_buffer(6612) := X"00000000";
		ram_buffer(6613) := X"00000000";
		ram_buffer(6614) := X"00000000";
		ram_buffer(6615) := X"00000000";
		ram_buffer(6616) := X"00000000";
		ram_buffer(6617) := X"00000000";
		ram_buffer(6618) := X"00000000";
		ram_buffer(6619) := X"00000000";
		ram_buffer(6620) := X"00000000";
		ram_buffer(6621) := X"00000000";
		ram_buffer(6622) := X"00000000";
		ram_buffer(6623) := X"00000000";
		ram_buffer(6624) := X"00000000";
		ram_buffer(6625) := X"00000000";
		ram_buffer(6626) := X"00000000";
		ram_buffer(6627) := X"00000000";
		ram_buffer(6628) := X"00000000";
		ram_buffer(6629) := X"00000000";
		ram_buffer(6630) := X"00000000";
		ram_buffer(6631) := X"00000000";
		ram_buffer(6632) := X"00000000";
		ram_buffer(6633) := X"00000000";
		ram_buffer(6634) := X"00000000";
		ram_buffer(6635) := X"00000000";
		ram_buffer(6636) := X"00000000";
		ram_buffer(6637) := X"00000000";
		ram_buffer(6638) := X"00000000";
		ram_buffer(6639) := X"00000000";
		ram_buffer(6640) := X"00000000";
		ram_buffer(6641) := X"00000000";
		ram_buffer(6642) := X"00000000";
		ram_buffer(6643) := X"00000000";
		ram_buffer(6644) := X"00000000";
		ram_buffer(6645) := X"00000000";
		ram_buffer(6646) := X"00000000";
		ram_buffer(6647) := X"00000000";
		ram_buffer(6648) := X"00000000";
		ram_buffer(6649) := X"00000000";
		ram_buffer(6650) := X"00000000";
		ram_buffer(6651) := X"00000000";
		ram_buffer(6652) := X"00000000";
		ram_buffer(6653) := X"00000000";
		ram_buffer(6654) := X"00000000";
		ram_buffer(6655) := X"00000000";
		ram_buffer(6656) := X"00000000";
		ram_buffer(6657) := X"00000000";
		ram_buffer(6658) := X"00000000";
		ram_buffer(6659) := X"00000000";
		ram_buffer(6660) := X"00000000";
		ram_buffer(6661) := X"00000000";
		ram_buffer(6662) := X"00000000";
		ram_buffer(6663) := X"00000000";
		ram_buffer(6664) := X"00000000";
		ram_buffer(6665) := X"00000000";
		ram_buffer(6666) := X"00000000";
		ram_buffer(6667) := X"00000000";
		ram_buffer(6668) := X"00000000";
		ram_buffer(6669) := X"00000000";
		ram_buffer(6670) := X"00000000";
		ram_buffer(6671) := X"00000000";
		ram_buffer(6672) := X"00000000";
		ram_buffer(6673) := X"00000000";
		ram_buffer(6674) := X"00000000";
		ram_buffer(6675) := X"00000000";
		ram_buffer(6676) := X"00000000";
		ram_buffer(6677) := X"00000000";
		ram_buffer(6678) := X"00000000";
		ram_buffer(6679) := X"00000000";
		ram_buffer(6680) := X"00000000";
		ram_buffer(6681) := X"00000000";
		ram_buffer(6682) := X"00000000";
		ram_buffer(6683) := X"00000000";
		ram_buffer(6684) := X"00000000";
		ram_buffer(6685) := X"00000000";
		ram_buffer(6686) := X"00000000";
		ram_buffer(6687) := X"00000000";
		ram_buffer(6688) := X"00000000";
		ram_buffer(6689) := X"00000000";
		ram_buffer(6690) := X"00000000";
		ram_buffer(6691) := X"00000000";
		ram_buffer(6692) := X"00000000";
		ram_buffer(6693) := X"00000000";
		ram_buffer(6694) := X"00000000";
		ram_buffer(6695) := X"00000000";
		ram_buffer(6696) := X"00000000";
		ram_buffer(6697) := X"00000000";
		ram_buffer(6698) := X"00000000";
		ram_buffer(6699) := X"00000000";
		ram_buffer(6700) := X"00000000";
		ram_buffer(6701) := X"00000000";
		ram_buffer(6702) := X"00000000";
		ram_buffer(6703) := X"00000000";
		ram_buffer(6704) := X"00000000";
		ram_buffer(6705) := X"00000000";
		ram_buffer(6706) := X"00000000";
		ram_buffer(6707) := X"00000000";
		ram_buffer(6708) := X"00000000";
		ram_buffer(6709) := X"00000000";
		ram_buffer(6710) := X"00000000";
		ram_buffer(6711) := X"00000000";
		ram_buffer(6712) := X"00000000";
		ram_buffer(6713) := X"00000000";
		ram_buffer(6714) := X"00000000";
		ram_buffer(6715) := X"00000000";
		ram_buffer(6716) := X"00000000";
		ram_buffer(6717) := X"00000000";
		ram_buffer(6718) := X"00000000";
		ram_buffer(6719) := X"00000000";
		ram_buffer(6720) := X"00000000";
		ram_buffer(6721) := X"00000000";
		ram_buffer(6722) := X"00000000";
		ram_buffer(6723) := X"00000000";
		ram_buffer(6724) := X"00000000";
		ram_buffer(6725) := X"00000000";
		ram_buffer(6726) := X"00000000";
		ram_buffer(6727) := X"00000000";
		ram_buffer(6728) := X"00000000";
		ram_buffer(6729) := X"00000000";
		ram_buffer(6730) := X"00000000";
		ram_buffer(6731) := X"00000000";
		ram_buffer(6732) := X"00000000";
		ram_buffer(6733) := X"00000000";
		ram_buffer(6734) := X"00000000";
		ram_buffer(6735) := X"00000000";
		ram_buffer(6736) := X"00000000";
		ram_buffer(6737) := X"00000000";
		ram_buffer(6738) := X"00000000";
		ram_buffer(6739) := X"00000000";
		ram_buffer(6740) := X"00000000";
		ram_buffer(6741) := X"00000000";
		ram_buffer(6742) := X"00000000";
		ram_buffer(6743) := X"00000000";
		ram_buffer(6744) := X"00000000";
		ram_buffer(6745) := X"00000000";
		ram_buffer(6746) := X"00000000";
		ram_buffer(6747) := X"00000000";
		ram_buffer(6748) := X"00000000";
		ram_buffer(6749) := X"00000000";
		ram_buffer(6750) := X"00000000";
		ram_buffer(6751) := X"00000000";
		ram_buffer(6752) := X"00000000";
		ram_buffer(6753) := X"00000000";
		ram_buffer(6754) := X"00000000";
		ram_buffer(6755) := X"00000000";
		ram_buffer(6756) := X"00000000";
		ram_buffer(6757) := X"00000000";
		ram_buffer(6758) := X"00000000";
		ram_buffer(6759) := X"00000000";
		ram_buffer(6760) := X"00000000";
		ram_buffer(6761) := X"00000000";
		ram_buffer(6762) := X"00000000";
		ram_buffer(6763) := X"00000000";
		ram_buffer(6764) := X"00000000";
		ram_buffer(6765) := X"00000000";
		ram_buffer(6766) := X"00000000";
		ram_buffer(6767) := X"00000000";
		ram_buffer(6768) := X"00000000";
		ram_buffer(6769) := X"00000000";
		ram_buffer(6770) := X"00000000";
		ram_buffer(6771) := X"00000000";
		ram_buffer(6772) := X"00000000";
		ram_buffer(6773) := X"00000000";
		ram_buffer(6774) := X"00000000";
		ram_buffer(6775) := X"00000000";
		ram_buffer(6776) := X"00000000";
		ram_buffer(6777) := X"00000000";
		ram_buffer(6778) := X"00000000";
		ram_buffer(6779) := X"00000000";
		ram_buffer(6780) := X"00000000";
		ram_buffer(6781) := X"00000000";
		ram_buffer(6782) := X"00000000";
		ram_buffer(6783) := X"00000000";
		ram_buffer(6784) := X"00000000";
		ram_buffer(6785) := X"00000000";
		ram_buffer(6786) := X"00000000";
		ram_buffer(6787) := X"00000000";
		ram_buffer(6788) := X"00000000";
		ram_buffer(6789) := X"00000000";
		ram_buffer(6790) := X"00000000";
		ram_buffer(6791) := X"00000000";
		ram_buffer(6792) := X"00000000";
		ram_buffer(6793) := X"00000000";
		ram_buffer(6794) := X"00000000";
		ram_buffer(6795) := X"00000000";
		ram_buffer(6796) := X"00000000";
		ram_buffer(6797) := X"00000000";
		ram_buffer(6798) := X"00000000";
		ram_buffer(6799) := X"00000000";
		ram_buffer(6800) := X"00000000";
		ram_buffer(6801) := X"00000000";
		ram_buffer(6802) := X"00000000";
		ram_buffer(6803) := X"00000000";
		ram_buffer(6804) := X"00000000";
		ram_buffer(6805) := X"00000000";
		ram_buffer(6806) := X"00000000";
		ram_buffer(6807) := X"00000000";
		ram_buffer(6808) := X"00000000";
		ram_buffer(6809) := X"00000000";
		ram_buffer(6810) := X"00000000";
		ram_buffer(6811) := X"00000000";
		ram_buffer(6812) := X"00000000";
		ram_buffer(6813) := X"00000000";
		ram_buffer(6814) := X"00000000";
		ram_buffer(6815) := X"00000000";
		ram_buffer(6816) := X"00000000";
		ram_buffer(6817) := X"00000000";
		ram_buffer(6818) := X"00000000";
		ram_buffer(6819) := X"00000000";
		ram_buffer(6820) := X"00000000";
		ram_buffer(6821) := X"00000000";
		ram_buffer(6822) := X"00000000";
		ram_buffer(6823) := X"00000000";
		ram_buffer(6824) := X"00000000";
		ram_buffer(6825) := X"00000000";
		ram_buffer(6826) := X"00000000";
		ram_buffer(6827) := X"00000000";
		ram_buffer(6828) := X"00000000";
		ram_buffer(6829) := X"00000000";
		ram_buffer(6830) := X"00000000";
		ram_buffer(6831) := X"00000000";
		ram_buffer(6832) := X"00000000";
		ram_buffer(6833) := X"00000000";
		ram_buffer(6834) := X"00000000";
		ram_buffer(6835) := X"00000000";
		ram_buffer(6836) := X"00000000";
		ram_buffer(6837) := X"00000000";
		ram_buffer(6838) := X"00000000";
		ram_buffer(6839) := X"00000000";
		ram_buffer(6840) := X"00000000";
		ram_buffer(6841) := X"00000000";
		ram_buffer(6842) := X"00000000";
		ram_buffer(6843) := X"00000000";
		ram_buffer(6844) := X"00000000";
		ram_buffer(6845) := X"00000000";
		ram_buffer(6846) := X"00000000";
		ram_buffer(6847) := X"00000000";
		ram_buffer(6848) := X"00000000";
		ram_buffer(6849) := X"00000000";
		ram_buffer(6850) := X"00000000";
		ram_buffer(6851) := X"00000000";
		ram_buffer(6852) := X"00000000";
		ram_buffer(6853) := X"00000000";
		ram_buffer(6854) := X"00000000";
		ram_buffer(6855) := X"00000000";
		ram_buffer(6856) := X"00000000";
		ram_buffer(6857) := X"00000000";
		ram_buffer(6858) := X"00000000";
		ram_buffer(6859) := X"00000000";
		ram_buffer(6860) := X"00000000";
		ram_buffer(6861) := X"00000000";
		ram_buffer(6862) := X"00000000";
		ram_buffer(6863) := X"00000000";
		ram_buffer(6864) := X"00000000";
		ram_buffer(6865) := X"00000000";
		ram_buffer(6866) := X"00000000";
		ram_buffer(6867) := X"00000000";
		ram_buffer(6868) := X"00000000";
		ram_buffer(6869) := X"00000000";
		ram_buffer(6870) := X"00000000";
		ram_buffer(6871) := X"00000000";
		ram_buffer(6872) := X"00000000";
		ram_buffer(6873) := X"00000000";
		ram_buffer(6874) := X"00000000";
		ram_buffer(6875) := X"00000000";
		ram_buffer(6876) := X"00000000";
		ram_buffer(6877) := X"00000000";
		ram_buffer(6878) := X"00000000";
		ram_buffer(6879) := X"00000000";
		ram_buffer(6880) := X"00000000";
		ram_buffer(6881) := X"00000000";
		ram_buffer(6882) := X"00000000";
		ram_buffer(6883) := X"00000000";
		ram_buffer(6884) := X"00000000";
		ram_buffer(6885) := X"00000000";
		ram_buffer(6886) := X"00000000";
		ram_buffer(6887) := X"00000000";
		ram_buffer(6888) := X"00000000";
		ram_buffer(6889) := X"00000000";
		ram_buffer(6890) := X"00000000";
		ram_buffer(6891) := X"00000000";
		ram_buffer(6892) := X"00000000";
		ram_buffer(6893) := X"00000000";
		ram_buffer(6894) := X"00000000";
		ram_buffer(6895) := X"00000000";
		ram_buffer(6896) := X"00000000";
		ram_buffer(6897) := X"00000000";
		ram_buffer(6898) := X"00000000";
		ram_buffer(6899) := X"00000000";
		ram_buffer(6900) := X"00000000";
		ram_buffer(6901) := X"00000000";
		ram_buffer(6902) := X"00000000";
		ram_buffer(6903) := X"00000000";
		ram_buffer(6904) := X"00000000";
		ram_buffer(6905) := X"00000000";
		ram_buffer(6906) := X"00000000";
		ram_buffer(6907) := X"00000000";
		ram_buffer(6908) := X"00000000";
		ram_buffer(6909) := X"00000000";
		ram_buffer(6910) := X"00000000";
		ram_buffer(6911) := X"00000000";
		ram_buffer(6912) := X"00000000";
		ram_buffer(6913) := X"00000000";
		ram_buffer(6914) := X"00000000";
		ram_buffer(6915) := X"00000000";
		ram_buffer(6916) := X"00000000";
		ram_buffer(6917) := X"00000000";
		ram_buffer(6918) := X"00000000";
		ram_buffer(6919) := X"00000000";
		ram_buffer(6920) := X"00000000";
		ram_buffer(6921) := X"00000000";
		ram_buffer(6922) := X"00000000";
		ram_buffer(6923) := X"00000000";
		ram_buffer(6924) := X"00000000";
		ram_buffer(6925) := X"00000000";
		ram_buffer(6926) := X"00000000";
		ram_buffer(6927) := X"00000000";
		ram_buffer(6928) := X"00000000";
		ram_buffer(6929) := X"00000000";
		ram_buffer(6930) := X"00000000";
		ram_buffer(6931) := X"00000000";
		ram_buffer(6932) := X"00000000";
		ram_buffer(6933) := X"00000000";
		ram_buffer(6934) := X"00000000";
		ram_buffer(6935) := X"00000000";
		ram_buffer(6936) := X"00000000";
		ram_buffer(6937) := X"00000000";
		ram_buffer(6938) := X"00000000";
		ram_buffer(6939) := X"00000000";
		ram_buffer(6940) := X"00000000";
		ram_buffer(6941) := X"00000000";
		ram_buffer(6942) := X"00000000";
		ram_buffer(6943) := X"00000000";
		ram_buffer(6944) := X"00000000";
		ram_buffer(6945) := X"00000000";
		ram_buffer(6946) := X"00000000";
		ram_buffer(6947) := X"00000000";
		ram_buffer(6948) := X"00000000";
		ram_buffer(6949) := X"00000000";
		ram_buffer(6950) := X"00000000";
		ram_buffer(6951) := X"00000000";
		ram_buffer(6952) := X"00000000";
		ram_buffer(6953) := X"00000000";
		ram_buffer(6954) := X"00000000";
		ram_buffer(6955) := X"00000000";
		ram_buffer(6956) := X"00000000";
		ram_buffer(6957) := X"00000000";
		ram_buffer(6958) := X"00000000";
		ram_buffer(6959) := X"00000000";
		ram_buffer(6960) := X"00000000";
		ram_buffer(6961) := X"00000000";
		ram_buffer(6962) := X"00000000";
		ram_buffer(6963) := X"00000000";
		ram_buffer(6964) := X"00000000";
		ram_buffer(6965) := X"00000000";
		ram_buffer(6966) := X"00000000";
		ram_buffer(6967) := X"00000000";
		ram_buffer(6968) := X"00000000";
		ram_buffer(6969) := X"00000000";
		ram_buffer(6970) := X"00000000";
		ram_buffer(6971) := X"00000000";
		ram_buffer(6972) := X"00000000";
		ram_buffer(6973) := X"00000000";
		ram_buffer(6974) := X"00000000";
		ram_buffer(6975) := X"00000000";
		ram_buffer(6976) := X"00000000";
		ram_buffer(6977) := X"00000000";
		ram_buffer(6978) := X"00000000";
		ram_buffer(6979) := X"00000000";
		ram_buffer(6980) := X"00000000";
		ram_buffer(6981) := X"00000000";
		ram_buffer(6982) := X"00000000";
		ram_buffer(6983) := X"00000000";
		ram_buffer(6984) := X"00000000";
		ram_buffer(6985) := X"00000000";
		ram_buffer(6986) := X"00000000";
		ram_buffer(6987) := X"00000000";
		ram_buffer(6988) := X"00000000";
		ram_buffer(6989) := X"00000000";
		ram_buffer(6990) := X"00000000";
		ram_buffer(6991) := X"00000000";
		ram_buffer(6992) := X"00000000";
		ram_buffer(6993) := X"00000000";
		ram_buffer(6994) := X"00000000";
		ram_buffer(6995) := X"00000000";
		ram_buffer(6996) := X"00000000";
		ram_buffer(6997) := X"00000000";
		ram_buffer(6998) := X"00000000";
		ram_buffer(6999) := X"00000000";
		ram_buffer(7000) := X"00000000";
		ram_buffer(7001) := X"00000000";
		ram_buffer(7002) := X"00000000";
		ram_buffer(7003) := X"00000000";
		ram_buffer(7004) := X"00000000";
		ram_buffer(7005) := X"00000000";
		ram_buffer(7006) := X"00000000";
		ram_buffer(7007) := X"00000000";
		ram_buffer(7008) := X"00000000";
		ram_buffer(7009) := X"00000000";
		ram_buffer(7010) := X"00000000";
		ram_buffer(7011) := X"00000000";
		ram_buffer(7012) := X"00000000";
		ram_buffer(7013) := X"00000000";
		ram_buffer(7014) := X"00000000";
		ram_buffer(7015) := X"00000000";
		ram_buffer(7016) := X"00000000";
		ram_buffer(7017) := X"00000000";
		ram_buffer(7018) := X"00000000";
		ram_buffer(7019) := X"00000000";
		ram_buffer(7020) := X"00000000";
		ram_buffer(7021) := X"00000000";
		ram_buffer(7022) := X"00000000";
		ram_buffer(7023) := X"00000000";
		ram_buffer(7024) := X"00000000";
		ram_buffer(7025) := X"00000000";
		ram_buffer(7026) := X"00000000";
		ram_buffer(7027) := X"00000000";
		ram_buffer(7028) := X"00000000";
		ram_buffer(7029) := X"00000000";
		ram_buffer(7030) := X"00000000";
		ram_buffer(7031) := X"00000000";
		ram_buffer(7032) := X"00000000";
		ram_buffer(7033) := X"00000000";
		ram_buffer(7034) := X"00000000";
		ram_buffer(7035) := X"00000000";
		ram_buffer(7036) := X"00000000";
		ram_buffer(7037) := X"00000000";
		ram_buffer(7038) := X"00000000";
		ram_buffer(7039) := X"00000000";
		ram_buffer(7040) := X"00000000";
		ram_buffer(7041) := X"00000000";
		ram_buffer(7042) := X"00000000";
		ram_buffer(7043) := X"00000000";
		ram_buffer(7044) := X"00000000";
		ram_buffer(7045) := X"00000000";
		ram_buffer(7046) := X"00000000";
		ram_buffer(7047) := X"00000000";
		ram_buffer(7048) := X"00000000";
		ram_buffer(7049) := X"00000000";
		ram_buffer(7050) := X"00000000";
		ram_buffer(7051) := X"00000000";
		ram_buffer(7052) := X"00000000";
		ram_buffer(7053) := X"00000000";
		ram_buffer(7054) := X"00000000";
		ram_buffer(7055) := X"00000000";
		ram_buffer(7056) := X"00000000";
		ram_buffer(7057) := X"00000000";
		ram_buffer(7058) := X"00000000";
		ram_buffer(7059) := X"00000000";
		ram_buffer(7060) := X"00000000";
		ram_buffer(7061) := X"00000000";
		ram_buffer(7062) := X"00000000";
		ram_buffer(7063) := X"00000000";
		ram_buffer(7064) := X"00000000";
		ram_buffer(7065) := X"00000000";
		ram_buffer(7066) := X"00000000";
		ram_buffer(7067) := X"00000000";
		ram_buffer(7068) := X"00000000";
		ram_buffer(7069) := X"00000000";
		ram_buffer(7070) := X"00000000";
		ram_buffer(7071) := X"00000000";
		ram_buffer(7072) := X"00000000";
		ram_buffer(7073) := X"00000000";
		ram_buffer(7074) := X"00000000";
		ram_buffer(7075) := X"00000000";
		ram_buffer(7076) := X"00000000";
		ram_buffer(7077) := X"00000000";
		ram_buffer(7078) := X"00000000";
		ram_buffer(7079) := X"00000000";
		ram_buffer(7080) := X"00000000";
		ram_buffer(7081) := X"00000000";
		ram_buffer(7082) := X"00000000";
		ram_buffer(7083) := X"00000000";
		ram_buffer(7084) := X"00000000";
		ram_buffer(7085) := X"00000000";
		ram_buffer(7086) := X"00000000";
		ram_buffer(7087) := X"00000000";
		ram_buffer(7088) := X"00000000";
		ram_buffer(7089) := X"00000000";
		ram_buffer(7090) := X"00000000";
		ram_buffer(7091) := X"00000000";
		ram_buffer(7092) := X"00000000";
		ram_buffer(7093) := X"00000000";
		ram_buffer(7094) := X"00000000";
		ram_buffer(7095) := X"00000000";
		ram_buffer(7096) := X"00000000";
		ram_buffer(7097) := X"00000000";
		ram_buffer(7098) := X"00000000";
		ram_buffer(7099) := X"00000000";
		ram_buffer(7100) := X"00000000";
		ram_buffer(7101) := X"00000000";
		ram_buffer(7102) := X"00000000";
		ram_buffer(7103) := X"00000000";
		ram_buffer(7104) := X"00000000";
		ram_buffer(7105) := X"00000000";
		ram_buffer(7106) := X"00000000";
		ram_buffer(7107) := X"00000000";
		ram_buffer(7108) := X"00000000";
		ram_buffer(7109) := X"00000000";
		ram_buffer(7110) := X"00000000";
		ram_buffer(7111) := X"00000000";
		ram_buffer(7112) := X"00000000";
		ram_buffer(7113) := X"00000000";
		ram_buffer(7114) := X"00000000";
		ram_buffer(7115) := X"00000000";
		ram_buffer(7116) := X"00000000";
		ram_buffer(7117) := X"00000000";
		ram_buffer(7118) := X"00000000";
		ram_buffer(7119) := X"00000000";
		ram_buffer(7120) := X"00000000";
		ram_buffer(7121) := X"00000000";
		ram_buffer(7122) := X"00000000";
		ram_buffer(7123) := X"00000000";
		ram_buffer(7124) := X"00000000";
		ram_buffer(7125) := X"00000000";
		ram_buffer(7126) := X"00000000";
		ram_buffer(7127) := X"00000000";
		ram_buffer(7128) := X"00000000";
		ram_buffer(7129) := X"00000000";
		ram_buffer(7130) := X"00000000";
		ram_buffer(7131) := X"00000000";
		ram_buffer(7132) := X"00000000";
		ram_buffer(7133) := X"00000000";
		ram_buffer(7134) := X"00000000";
		ram_buffer(7135) := X"00000000";
		ram_buffer(7136) := X"00000000";
		ram_buffer(7137) := X"00000000";
		ram_buffer(7138) := X"00000000";
		ram_buffer(7139) := X"00000000";
		ram_buffer(7140) := X"00000000";
		ram_buffer(7141) := X"00000000";
		ram_buffer(7142) := X"00000000";
		ram_buffer(7143) := X"00000000";
		ram_buffer(7144) := X"00000000";
		ram_buffer(7145) := X"00000000";
		ram_buffer(7146) := X"00000000";
		ram_buffer(7147) := X"00000000";
		ram_buffer(7148) := X"00000000";
		ram_buffer(7149) := X"00000000";
		ram_buffer(7150) := X"00000000";
		ram_buffer(7151) := X"00000000";
		ram_buffer(7152) := X"00000000";
		ram_buffer(7153) := X"00000000";
		ram_buffer(7154) := X"00000000";
		ram_buffer(7155) := X"00000000";
		ram_buffer(7156) := X"00000000";
		ram_buffer(7157) := X"00000000";
		ram_buffer(7158) := X"00000000";
		ram_buffer(7159) := X"00000000";
		ram_buffer(7160) := X"00000000";
		ram_buffer(7161) := X"00000000";
		ram_buffer(7162) := X"00000000";
		ram_buffer(7163) := X"00000000";
		ram_buffer(7164) := X"00000000";
		ram_buffer(7165) := X"00000000";
		ram_buffer(7166) := X"00000000";
		ram_buffer(7167) := X"00000000";
		ram_buffer(7168) := X"00000000";
		ram_buffer(7169) := X"00000000";
		ram_buffer(7170) := X"00000000";
		ram_buffer(7171) := X"00000000";
		ram_buffer(7172) := X"00000000";
		ram_buffer(7173) := X"00000000";
		ram_buffer(7174) := X"00000000";
		ram_buffer(7175) := X"00000000";
		ram_buffer(7176) := X"00000000";
		ram_buffer(7177) := X"00000000";
		ram_buffer(7178) := X"00000000";
		ram_buffer(7179) := X"00000000";
		ram_buffer(7180) := X"00000000";
		ram_buffer(7181) := X"00000000";
		ram_buffer(7182) := X"00000000";
		ram_buffer(7183) := X"00000000";
		ram_buffer(7184) := X"00000000";
		ram_buffer(7185) := X"00000000";
		ram_buffer(7186) := X"00000000";
		ram_buffer(7187) := X"00000000";
		ram_buffer(7188) := X"00000000";
		ram_buffer(7189) := X"00000000";
		ram_buffer(7190) := X"00000000";
		ram_buffer(7191) := X"00000000";
		ram_buffer(7192) := X"00000000";
		ram_buffer(7193) := X"00000000";
		ram_buffer(7194) := X"00000000";
		ram_buffer(7195) := X"00000000";
		ram_buffer(7196) := X"00000000";
		ram_buffer(7197) := X"00000000";
		ram_buffer(7198) := X"00000000";
		ram_buffer(7199) := X"00000000";
		ram_buffer(7200) := X"00000000";
		ram_buffer(7201) := X"00000000";
		ram_buffer(7202) := X"00000000";
		ram_buffer(7203) := X"00000000";
		ram_buffer(7204) := X"00000000";
		ram_buffer(7205) := X"00000000";
		ram_buffer(7206) := X"00000000";
		ram_buffer(7207) := X"00000000";
		ram_buffer(7208) := X"00000000";
		ram_buffer(7209) := X"00000000";
		ram_buffer(7210) := X"00000000";
		ram_buffer(7211) := X"00000000";
		ram_buffer(7212) := X"00000000";
		ram_buffer(7213) := X"00000000";
		ram_buffer(7214) := X"00000000";
		ram_buffer(7215) := X"00000000";
		ram_buffer(7216) := X"00000000";
		ram_buffer(7217) := X"00000000";
		ram_buffer(7218) := X"00000000";
		ram_buffer(7219) := X"00000000";
		ram_buffer(7220) := X"00000000";
		ram_buffer(7221) := X"00000000";
		ram_buffer(7222) := X"00000000";
		ram_buffer(7223) := X"00000000";
		ram_buffer(7224) := X"00000000";
		ram_buffer(7225) := X"00000000";
		ram_buffer(7226) := X"00000000";
		ram_buffer(7227) := X"00000000";
		ram_buffer(7228) := X"00000000";
		ram_buffer(7229) := X"00000000";
		ram_buffer(7230) := X"00000000";
		ram_buffer(7231) := X"00000000";
		ram_buffer(7232) := X"00000000";
		ram_buffer(7233) := X"00000000";
		ram_buffer(7234) := X"00000000";
		ram_buffer(7235) := X"00000000";
		ram_buffer(7236) := X"00000000";
		ram_buffer(7237) := X"00000000";
		ram_buffer(7238) := X"00000000";
		ram_buffer(7239) := X"00000000";
		ram_buffer(7240) := X"00000000";
		ram_buffer(7241) := X"00000000";
		ram_buffer(7242) := X"00000000";
		ram_buffer(7243) := X"00000000";
		ram_buffer(7244) := X"00000000";
		ram_buffer(7245) := X"00000000";
		ram_buffer(7246) := X"00000000";
		ram_buffer(7247) := X"00000000";
		ram_buffer(7248) := X"00000000";
		ram_buffer(7249) := X"00000000";
		ram_buffer(7250) := X"00000000";
		ram_buffer(7251) := X"00000000";
		ram_buffer(7252) := X"00000000";
		ram_buffer(7253) := X"00000000";
		ram_buffer(7254) := X"00000000";
		ram_buffer(7255) := X"00000000";
		ram_buffer(7256) := X"00000000";
		ram_buffer(7257) := X"00000000";
		ram_buffer(7258) := X"00000000";
		ram_buffer(7259) := X"00000000";
		ram_buffer(7260) := X"00000000";
		ram_buffer(7261) := X"00000000";
		ram_buffer(7262) := X"00000000";
		ram_buffer(7263) := X"00000000";
		ram_buffer(7264) := X"00000000";
		ram_buffer(7265) := X"00000000";
		ram_buffer(7266) := X"00000000";
		ram_buffer(7267) := X"00000000";
		ram_buffer(7268) := X"00000000";
		ram_buffer(7269) := X"00000000";
		ram_buffer(7270) := X"00000000";
		ram_buffer(7271) := X"00000000";
		ram_buffer(7272) := X"00000000";
		ram_buffer(7273) := X"00000000";
		ram_buffer(7274) := X"00000000";
		ram_buffer(7275) := X"00000000";
		ram_buffer(7276) := X"00000000";
		ram_buffer(7277) := X"00000000";
		ram_buffer(7278) := X"00000000";
		ram_buffer(7279) := X"00000000";
		ram_buffer(7280) := X"00000000";
		ram_buffer(7281) := X"00000000";
		ram_buffer(7282) := X"00000000";
		ram_buffer(7283) := X"00000000";
		ram_buffer(7284) := X"00000000";
		ram_buffer(7285) := X"00000000";
		ram_buffer(7286) := X"00000000";
		ram_buffer(7287) := X"00000000";
		ram_buffer(7288) := X"00000000";
		ram_buffer(7289) := X"00000000";
		ram_buffer(7290) := X"00000000";
		ram_buffer(7291) := X"00000000";
		ram_buffer(7292) := X"00000000";
		ram_buffer(7293) := X"00000000";
		ram_buffer(7294) := X"00000000";
		ram_buffer(7295) := X"00000000";
		ram_buffer(7296) := X"00000000";
		ram_buffer(7297) := X"00000000";
		ram_buffer(7298) := X"00000000";
		ram_buffer(7299) := X"00000000";
		ram_buffer(7300) := X"00000000";
		ram_buffer(7301) := X"00000000";
		ram_buffer(7302) := X"00000000";
		ram_buffer(7303) := X"00000000";
		ram_buffer(7304) := X"00000000";
		ram_buffer(7305) := X"00000000";
		ram_buffer(7306) := X"00000000";
		ram_buffer(7307) := X"00000000";
		ram_buffer(7308) := X"00000000";
		ram_buffer(7309) := X"00000000";
		ram_buffer(7310) := X"00000000";
		ram_buffer(7311) := X"00000000";
		ram_buffer(7312) := X"00000000";
		ram_buffer(7313) := X"00000000";
		ram_buffer(7314) := X"00000000";
		ram_buffer(7315) := X"00000000";
		ram_buffer(7316) := X"00000000";
		ram_buffer(7317) := X"00000000";
		ram_buffer(7318) := X"00000000";
		ram_buffer(7319) := X"00000000";
		ram_buffer(7320) := X"00000000";
		ram_buffer(7321) := X"00000000";
		ram_buffer(7322) := X"00000000";
		ram_buffer(7323) := X"00000000";
		ram_buffer(7324) := X"00000000";
		ram_buffer(7325) := X"00000000";
		ram_buffer(7326) := X"00000000";
		ram_buffer(7327) := X"00000000";
		ram_buffer(7328) := X"00000000";
		ram_buffer(7329) := X"00000000";
		ram_buffer(7330) := X"00000000";
		ram_buffer(7331) := X"00000000";
		ram_buffer(7332) := X"00000000";
		ram_buffer(7333) := X"00000000";
		ram_buffer(7334) := X"00000000";
		ram_buffer(7335) := X"00000000";
		ram_buffer(7336) := X"00000000";
		ram_buffer(7337) := X"00000000";
		ram_buffer(7338) := X"00000000";
		ram_buffer(7339) := X"00000000";
		ram_buffer(7340) := X"00000000";
		ram_buffer(7341) := X"00000000";
		ram_buffer(7342) := X"00000000";
		ram_buffer(7343) := X"00000000";
		ram_buffer(7344) := X"00000000";
		ram_buffer(7345) := X"00000000";
		ram_buffer(7346) := X"00000000";
		ram_buffer(7347) := X"00000000";
		ram_buffer(7348) := X"00000000";
		ram_buffer(7349) := X"00000000";
		ram_buffer(7350) := X"00000000";
		ram_buffer(7351) := X"00000000";
		ram_buffer(7352) := X"00000000";
		ram_buffer(7353) := X"00000000";
		ram_buffer(7354) := X"00000000";
		ram_buffer(7355) := X"00000000";
		ram_buffer(7356) := X"00000000";
		ram_buffer(7357) := X"00000000";
		ram_buffer(7358) := X"00000000";
		ram_buffer(7359) := X"00000000";
		ram_buffer(7360) := X"00000000";
		ram_buffer(7361) := X"00000000";
		ram_buffer(7362) := X"00000000";
		ram_buffer(7363) := X"00000000";
		ram_buffer(7364) := X"00000000";
		ram_buffer(7365) := X"00000000";
		ram_buffer(7366) := X"00000000";
		ram_buffer(7367) := X"00000000";
		ram_buffer(7368) := X"00000000";
		ram_buffer(7369) := X"00000000";
		ram_buffer(7370) := X"00000000";
		ram_buffer(7371) := X"00000000";
		ram_buffer(7372) := X"00000000";
		ram_buffer(7373) := X"00000000";
		ram_buffer(7374) := X"00000000";
		ram_buffer(7375) := X"00000000";
		ram_buffer(7376) := X"00000000";
		ram_buffer(7377) := X"00000000";
		ram_buffer(7378) := X"00000000";
		ram_buffer(7379) := X"00000000";
		ram_buffer(7380) := X"00000000";
		ram_buffer(7381) := X"00000000";
		ram_buffer(7382) := X"00000000";
		ram_buffer(7383) := X"00000000";
		ram_buffer(7384) := X"00000000";
		ram_buffer(7385) := X"00000000";
		ram_buffer(7386) := X"00000000";
		ram_buffer(7387) := X"00000000";
		ram_buffer(7388) := X"00000000";
		ram_buffer(7389) := X"00000000";
		ram_buffer(7390) := X"00000000";
		ram_buffer(7391) := X"00000000";
		ram_buffer(7392) := X"00000000";
		ram_buffer(7393) := X"00000000";
		ram_buffer(7394) := X"00000000";
		ram_buffer(7395) := X"00000000";
		ram_buffer(7396) := X"00000000";
		ram_buffer(7397) := X"00000000";
		ram_buffer(7398) := X"00000000";
		ram_buffer(7399) := X"00000000";
		ram_buffer(7400) := X"00000000";
		ram_buffer(7401) := X"00000000";
		ram_buffer(7402) := X"00000000";
		ram_buffer(7403) := X"00000000";
		ram_buffer(7404) := X"00000000";
		ram_buffer(7405) := X"00000000";
		ram_buffer(7406) := X"00000000";
		ram_buffer(7407) := X"00000000";
		ram_buffer(7408) := X"00000000";
		ram_buffer(7409) := X"00000000";
		ram_buffer(7410) := X"00000000";
		ram_buffer(7411) := X"00000000";
		ram_buffer(7412) := X"00000000";
		ram_buffer(7413) := X"00000000";
		ram_buffer(7414) := X"00000000";
		ram_buffer(7415) := X"00000000";
		ram_buffer(7416) := X"00000000";
		ram_buffer(7417) := X"00000000";
		ram_buffer(7418) := X"00000000";
		ram_buffer(7419) := X"00000000";
		ram_buffer(7420) := X"00000000";
		ram_buffer(7421) := X"00000000";
		ram_buffer(7422) := X"00000000";
		ram_buffer(7423) := X"00000000";
		ram_buffer(7424) := X"00000000";
		ram_buffer(7425) := X"00000000";
		ram_buffer(7426) := X"00000000";
		ram_buffer(7427) := X"00000000";
		ram_buffer(7428) := X"00000000";
		ram_buffer(7429) := X"00000000";
		ram_buffer(7430) := X"00000000";
		ram_buffer(7431) := X"00000000";
		ram_buffer(7432) := X"00000000";
		ram_buffer(7433) := X"00000000";
		ram_buffer(7434) := X"00000000";
		ram_buffer(7435) := X"00000000";
		ram_buffer(7436) := X"00000000";
		ram_buffer(7437) := X"00000000";
		ram_buffer(7438) := X"00000000";
		ram_buffer(7439) := X"00000000";
		ram_buffer(7440) := X"00000000";
		ram_buffer(7441) := X"00000000";
		ram_buffer(7442) := X"00000000";
		ram_buffer(7443) := X"00000000";
		ram_buffer(7444) := X"00000000";
		ram_buffer(7445) := X"00000000";
		ram_buffer(7446) := X"00000000";
		ram_buffer(7447) := X"00000000";
		ram_buffer(7448) := X"00000000";
		ram_buffer(7449) := X"00000000";
		ram_buffer(7450) := X"00000000";
		ram_buffer(7451) := X"00000000";
		ram_buffer(7452) := X"00000000";
		ram_buffer(7453) := X"00000000";
		ram_buffer(7454) := X"00000000";
		ram_buffer(7455) := X"00000000";
		ram_buffer(7456) := X"00000000";
		ram_buffer(7457) := X"00000000";
		ram_buffer(7458) := X"00000000";
		ram_buffer(7459) := X"00000000";
		ram_buffer(7460) := X"00000000";
		ram_buffer(7461) := X"00000000";
		ram_buffer(7462) := X"00000000";
		ram_buffer(7463) := X"00000000";
		ram_buffer(7464) := X"00000000";
		ram_buffer(7465) := X"00000000";
		ram_buffer(7466) := X"00000000";
		ram_buffer(7467) := X"00000000";
		ram_buffer(7468) := X"00000000";
		ram_buffer(7469) := X"00000000";
		ram_buffer(7470) := X"00000000";
		ram_buffer(7471) := X"00000000";
		ram_buffer(7472) := X"00000000";
		ram_buffer(7473) := X"00000000";
		ram_buffer(7474) := X"00000000";
		ram_buffer(7475) := X"00000000";
		ram_buffer(7476) := X"00000000";
		ram_buffer(7477) := X"00000000";
		ram_buffer(7478) := X"00000000";
		ram_buffer(7479) := X"00000000";
		ram_buffer(7480) := X"00000000";
		ram_buffer(7481) := X"00000000";
		ram_buffer(7482) := X"00000000";
		ram_buffer(7483) := X"00000000";
		ram_buffer(7484) := X"00000000";
		ram_buffer(7485) := X"00000000";
		ram_buffer(7486) := X"00000000";
		ram_buffer(7487) := X"00000000";
		ram_buffer(7488) := X"00000000";
		ram_buffer(7489) := X"00000000";
		ram_buffer(7490) := X"00000000";
		ram_buffer(7491) := X"00000000";
		ram_buffer(7492) := X"00000000";
		ram_buffer(7493) := X"00000000";
		ram_buffer(7494) := X"00000000";
		ram_buffer(7495) := X"00000000";
		ram_buffer(7496) := X"00000000";
		ram_buffer(7497) := X"00000000";
		ram_buffer(7498) := X"00000000";
		ram_buffer(7499) := X"00000000";
		ram_buffer(7500) := X"00000000";
		ram_buffer(7501) := X"00000000";
		ram_buffer(7502) := X"00000000";
		ram_buffer(7503) := X"00000000";
		ram_buffer(7504) := X"00000000";
		ram_buffer(7505) := X"00000000";
		ram_buffer(7506) := X"00000000";
		ram_buffer(7507) := X"00000000";
		ram_buffer(7508) := X"00000000";
		ram_buffer(7509) := X"00000000";
		ram_buffer(7510) := X"00000000";
		ram_buffer(7511) := X"00000000";
		ram_buffer(7512) := X"00000000";
		ram_buffer(7513) := X"00000000";
		ram_buffer(7514) := X"00000000";
		ram_buffer(7515) := X"00000000";
		ram_buffer(7516) := X"00000000";
		ram_buffer(7517) := X"00000000";
		ram_buffer(7518) := X"00000000";
		ram_buffer(7519) := X"00000000";
		ram_buffer(7520) := X"00000000";
		ram_buffer(7521) := X"00000000";
		ram_buffer(7522) := X"00000000";
		ram_buffer(7523) := X"00000000";
		ram_buffer(7524) := X"00000000";
		ram_buffer(7525) := X"00000000";
		ram_buffer(7526) := X"00000000";
		ram_buffer(7527) := X"00000000";
		ram_buffer(7528) := X"00000000";
		ram_buffer(7529) := X"00000000";
		ram_buffer(7530) := X"00000000";
		ram_buffer(7531) := X"00000000";
		ram_buffer(7532) := X"00000000";
		ram_buffer(7533) := X"00000000";
		ram_buffer(7534) := X"00000000";
		ram_buffer(7535) := X"00000000";
		ram_buffer(7536) := X"00000000";
		ram_buffer(7537) := X"00000000";
		ram_buffer(7538) := X"00000000";
		ram_buffer(7539) := X"00000000";
		ram_buffer(7540) := X"00000000";
		ram_buffer(7541) := X"00000000";
		ram_buffer(7542) := X"00000000";
		ram_buffer(7543) := X"00000000";
		ram_buffer(7544) := X"00000000";
		ram_buffer(7545) := X"00000000";
		ram_buffer(7546) := X"00000000";
		ram_buffer(7547) := X"00000000";
		ram_buffer(7548) := X"00000000";
		ram_buffer(7549) := X"00000000";
		ram_buffer(7550) := X"00000000";
		ram_buffer(7551) := X"00000000";
		ram_buffer(7552) := X"00000000";
		ram_buffer(7553) := X"00000000";
		ram_buffer(7554) := X"00000000";
		ram_buffer(7555) := X"00000000";
		ram_buffer(7556) := X"00000000";
		ram_buffer(7557) := X"00000000";
		ram_buffer(7558) := X"00000000";
		ram_buffer(7559) := X"00000000";
		ram_buffer(7560) := X"00000000";
		ram_buffer(7561) := X"00000000";
		ram_buffer(7562) := X"00000000";
		ram_buffer(7563) := X"00000000";
		ram_buffer(7564) := X"00000000";
		ram_buffer(7565) := X"00000000";
		ram_buffer(7566) := X"00000000";
		ram_buffer(7567) := X"00000000";
		ram_buffer(7568) := X"00000000";
		ram_buffer(7569) := X"00000000";
		ram_buffer(7570) := X"00000000";
		ram_buffer(7571) := X"00000000";
		ram_buffer(7572) := X"00000000";
		ram_buffer(7573) := X"00000000";
		ram_buffer(7574) := X"00000000";
		ram_buffer(7575) := X"00000000";
		ram_buffer(7576) := X"00000000";
		ram_buffer(7577) := X"00000000";
		ram_buffer(7578) := X"00000000";
		ram_buffer(7579) := X"00000000";
		ram_buffer(7580) := X"00000000";
		ram_buffer(7581) := X"00000000";
		ram_buffer(7582) := X"00000000";
		ram_buffer(7583) := X"00000000";
		ram_buffer(7584) := X"00000000";
		ram_buffer(7585) := X"00000000";
		ram_buffer(7586) := X"00000000";
		ram_buffer(7587) := X"00000000";
		ram_buffer(7588) := X"00000000";
		ram_buffer(7589) := X"00000000";
		ram_buffer(7590) := X"00000000";
		ram_buffer(7591) := X"00000000";
		ram_buffer(7592) := X"00000000";
		ram_buffer(7593) := X"00000000";
		ram_buffer(7594) := X"00000000";
		ram_buffer(7595) := X"00000000";
		ram_buffer(7596) := X"00000000";
		ram_buffer(7597) := X"00000000";
		ram_buffer(7598) := X"00000000";
		ram_buffer(7599) := X"00000000";
		ram_buffer(7600) := X"00000000";
		ram_buffer(7601) := X"00000000";
		ram_buffer(7602) := X"00000000";
		ram_buffer(7603) := X"00000000";
		ram_buffer(7604) := X"00000000";
		ram_buffer(7605) := X"00000000";
		ram_buffer(7606) := X"00000000";
		ram_buffer(7607) := X"00000000";
		ram_buffer(7608) := X"00000000";
		ram_buffer(7609) := X"00000000";
		ram_buffer(7610) := X"00000000";
		ram_buffer(7611) := X"00000000";
		ram_buffer(7612) := X"00000000";
		ram_buffer(7613) := X"00000000";
		ram_buffer(7614) := X"00000000";
		ram_buffer(7615) := X"00000000";
		ram_buffer(7616) := X"00000000";
		ram_buffer(7617) := X"00000000";
		ram_buffer(7618) := X"00000000";
		ram_buffer(7619) := X"00000000";
		ram_buffer(7620) := X"00000000";
		ram_buffer(7621) := X"00000000";
		ram_buffer(7622) := X"00000000";
		ram_buffer(7623) := X"00000000";
		ram_buffer(7624) := X"00000000";
		ram_buffer(7625) := X"00000000";
		ram_buffer(7626) := X"00000000";
		ram_buffer(7627) := X"00000000";
		ram_buffer(7628) := X"00000000";
		ram_buffer(7629) := X"00000000";
		ram_buffer(7630) := X"00000000";
		ram_buffer(7631) := X"00000000";
		ram_buffer(7632) := X"00000000";
		ram_buffer(7633) := X"00000000";
		ram_buffer(7634) := X"00000000";
		ram_buffer(7635) := X"00000000";
		ram_buffer(7636) := X"00000000";
		ram_buffer(7637) := X"00000000";
		ram_buffer(7638) := X"00000000";
		ram_buffer(7639) := X"00000000";
		ram_buffer(7640) := X"00000000";
		ram_buffer(7641) := X"00000000";
		ram_buffer(7642) := X"00000000";
		ram_buffer(7643) := X"00000000";
		ram_buffer(7644) := X"00000000";
		ram_buffer(7645) := X"00000000";
		ram_buffer(7646) := X"00000000";
		ram_buffer(7647) := X"00000000";
		ram_buffer(7648) := X"00000000";
		ram_buffer(7649) := X"00000000";
		ram_buffer(7650) := X"00000000";
		ram_buffer(7651) := X"00000000";
		ram_buffer(7652) := X"00000000";
		ram_buffer(7653) := X"00000000";
		ram_buffer(7654) := X"00000000";
		ram_buffer(7655) := X"00000000";
		ram_buffer(7656) := X"00000000";
		ram_buffer(7657) := X"00000000";
		ram_buffer(7658) := X"00000000";
		ram_buffer(7659) := X"00000000";
		ram_buffer(7660) := X"00000000";
		ram_buffer(7661) := X"00000000";
		ram_buffer(7662) := X"00000000";
		ram_buffer(7663) := X"00000000";
		ram_buffer(7664) := X"00000000";
		ram_buffer(7665) := X"00000000";
		ram_buffer(7666) := X"00000000";
		ram_buffer(7667) := X"00000000";
		ram_buffer(7668) := X"00000000";
		ram_buffer(7669) := X"00000000";
		ram_buffer(7670) := X"00000000";
		ram_buffer(7671) := X"00000000";
		ram_buffer(7672) := X"00000000";
		ram_buffer(7673) := X"00000000";
		ram_buffer(7674) := X"00000000";
		ram_buffer(7675) := X"00000000";
		ram_buffer(7676) := X"00000000";
		ram_buffer(7677) := X"00000000";
		ram_buffer(7678) := X"00000000";
		ram_buffer(7679) := X"00000000";
		ram_buffer(7680) := X"00000000";
		ram_buffer(7681) := X"00000000";
		ram_buffer(7682) := X"00000000";
		ram_buffer(7683) := X"00000000";
		ram_buffer(7684) := X"00000000";
		ram_buffer(7685) := X"00000000";
		ram_buffer(7686) := X"00000000";
		ram_buffer(7687) := X"00000000";
		ram_buffer(7688) := X"00000000";
		ram_buffer(7689) := X"00000000";
		ram_buffer(7690) := X"00000000";
		ram_buffer(7691) := X"00000000";
		ram_buffer(7692) := X"00000000";
		ram_buffer(7693) := X"00000000";
		ram_buffer(7694) := X"00000000";
		ram_buffer(7695) := X"00000000";
		ram_buffer(7696) := X"00000000";
		ram_buffer(7697) := X"00000000";
		ram_buffer(7698) := X"00000000";
		ram_buffer(7699) := X"00000000";
		ram_buffer(7700) := X"00000000";
		ram_buffer(7701) := X"00000000";
		ram_buffer(7702) := X"00000000";
		ram_buffer(7703) := X"00000000";
		ram_buffer(7704) := X"00000000";
		ram_buffer(7705) := X"00000000";
		ram_buffer(7706) := X"00000000";
		ram_buffer(7707) := X"00000000";
		ram_buffer(7708) := X"00000000";
		ram_buffer(7709) := X"00000000";
		ram_buffer(7710) := X"00000000";
		ram_buffer(7711) := X"00000000";
		ram_buffer(7712) := X"00000000";
		ram_buffer(7713) := X"00000000";
		ram_buffer(7714) := X"00000000";
		ram_buffer(7715) := X"00000000";
		ram_buffer(7716) := X"00000000";
		ram_buffer(7717) := X"00000000";
		ram_buffer(7718) := X"00000000";
		ram_buffer(7719) := X"00000000";
		ram_buffer(7720) := X"00000000";
		ram_buffer(7721) := X"00000000";
		ram_buffer(7722) := X"00000000";
		ram_buffer(7723) := X"00000000";
		ram_buffer(7724) := X"00000000";
		ram_buffer(7725) := X"00000000";
		ram_buffer(7726) := X"00000000";
		ram_buffer(7727) := X"00000000";
		ram_buffer(7728) := X"00000000";
		ram_buffer(7729) := X"00000000";
		ram_buffer(7730) := X"00000000";
		ram_buffer(7731) := X"00000000";
		ram_buffer(7732) := X"00000000";
		ram_buffer(7733) := X"00000000";
		ram_buffer(7734) := X"00000000";
		ram_buffer(7735) := X"00000000";
		ram_buffer(7736) := X"00000000";
		ram_buffer(7737) := X"00000000";
		ram_buffer(7738) := X"00000000";
		ram_buffer(7739) := X"00000000";
		ram_buffer(7740) := X"00000000";
		ram_buffer(7741) := X"00000000";
		ram_buffer(7742) := X"00000000";
		ram_buffer(7743) := X"00000000";
		ram_buffer(7744) := X"00000000";
		ram_buffer(7745) := X"00000000";
		ram_buffer(7746) := X"00000000";
		ram_buffer(7747) := X"00000000";
		ram_buffer(7748) := X"00000000";
		ram_buffer(7749) := X"00000000";
		ram_buffer(7750) := X"00000000";
		ram_buffer(7751) := X"00000000";
		ram_buffer(7752) := X"00000000";
		ram_buffer(7753) := X"00000000";
		ram_buffer(7754) := X"00000000";
		ram_buffer(7755) := X"00000000";
		ram_buffer(7756) := X"00000000";
		ram_buffer(7757) := X"00000000";
		ram_buffer(7758) := X"00000000";
		ram_buffer(7759) := X"00000000";
		ram_buffer(7760) := X"00000000";
		ram_buffer(7761) := X"00000000";
		ram_buffer(7762) := X"00000000";
		ram_buffer(7763) := X"00000000";
		ram_buffer(7764) := X"00000000";
		ram_buffer(7765) := X"00000000";
		ram_buffer(7766) := X"00000000";
		ram_buffer(7767) := X"00000000";
		ram_buffer(7768) := X"00000000";
		ram_buffer(7769) := X"00000000";
		ram_buffer(7770) := X"00000000";
		ram_buffer(7771) := X"00000000";
		ram_buffer(7772) := X"00000000";
		ram_buffer(7773) := X"00000000";
		ram_buffer(7774) := X"00000000";
		ram_buffer(7775) := X"00000000";
		ram_buffer(7776) := X"00000000";
		ram_buffer(7777) := X"00000000";
		ram_buffer(7778) := X"00000000";
		ram_buffer(7779) := X"00000000";
		ram_buffer(7780) := X"00000000";
		ram_buffer(7781) := X"00000000";
		ram_buffer(7782) := X"00000000";
		ram_buffer(7783) := X"00000000";
		ram_buffer(7784) := X"00000000";
		ram_buffer(7785) := X"00000000";
		ram_buffer(7786) := X"00000000";
		ram_buffer(7787) := X"00000000";
		ram_buffer(7788) := X"00000000";
		ram_buffer(7789) := X"00000000";
		ram_buffer(7790) := X"00000000";
		ram_buffer(7791) := X"00000000";
		ram_buffer(7792) := X"00000000";
		ram_buffer(7793) := X"00000000";
		ram_buffer(7794) := X"00000000";
		ram_buffer(7795) := X"00000000";
		ram_buffer(7796) := X"00000000";
		ram_buffer(7797) := X"00000000";
		ram_buffer(7798) := X"00000000";
		ram_buffer(7799) := X"00000000";
		ram_buffer(7800) := X"00000000";
		ram_buffer(7801) := X"00000000";
		ram_buffer(7802) := X"00000000";
		ram_buffer(7803) := X"00000000";
		ram_buffer(7804) := X"00000000";
		ram_buffer(7805) := X"00000000";
		ram_buffer(7806) := X"00000000";
		ram_buffer(7807) := X"00000000";
		ram_buffer(7808) := X"00000000";
		ram_buffer(7809) := X"00000000";
		ram_buffer(7810) := X"00000000";
		ram_buffer(7811) := X"00000000";
		ram_buffer(7812) := X"00000000";
		ram_buffer(7813) := X"00000000";
		ram_buffer(7814) := X"00000000";
		ram_buffer(7815) := X"00000000";
		ram_buffer(7816) := X"00000000";
		ram_buffer(7817) := X"00000000";
		ram_buffer(7818) := X"00000000";
		ram_buffer(7819) := X"00000000";
		ram_buffer(7820) := X"00000000";
		ram_buffer(7821) := X"00000000";
		ram_buffer(7822) := X"00000000";
		ram_buffer(7823) := X"00000000";
		ram_buffer(7824) := X"00000000";
		ram_buffer(7825) := X"00000000";
		ram_buffer(7826) := X"00000000";
		ram_buffer(7827) := X"00000000";
		ram_buffer(7828) := X"00000000";
		ram_buffer(7829) := X"00000000";
		ram_buffer(7830) := X"00000000";
		ram_buffer(7831) := X"00000000";
		ram_buffer(7832) := X"00000000";
		ram_buffer(7833) := X"00000000";
		ram_buffer(7834) := X"00000000";
		ram_buffer(7835) := X"00000000";
		ram_buffer(7836) := X"00000000";
		ram_buffer(7837) := X"00000000";
		ram_buffer(7838) := X"00000000";
		ram_buffer(7839) := X"00000000";
		ram_buffer(7840) := X"00000000";
		ram_buffer(7841) := X"00000000";
		ram_buffer(7842) := X"00000000";
		ram_buffer(7843) := X"00000000";
		ram_buffer(7844) := X"00000000";
		ram_buffer(7845) := X"00000000";
		ram_buffer(7846) := X"00000000";
		ram_buffer(7847) := X"00000000";
		ram_buffer(7848) := X"00000000";
		ram_buffer(7849) := X"00000000";
		ram_buffer(7850) := X"00000000";
		ram_buffer(7851) := X"00000000";
		ram_buffer(7852) := X"00000000";
		ram_buffer(7853) := X"00000000";
		ram_buffer(7854) := X"00000000";
		ram_buffer(7855) := X"00000000";
		ram_buffer(7856) := X"00000000";
		ram_buffer(7857) := X"00000000";
		ram_buffer(7858) := X"00000000";
		ram_buffer(7859) := X"00000000";
		ram_buffer(7860) := X"00000000";
		ram_buffer(7861) := X"00000000";
		ram_buffer(7862) := X"00000000";
		ram_buffer(7863) := X"00000000";
		ram_buffer(7864) := X"00000000";
		ram_buffer(7865) := X"00000000";
		ram_buffer(7866) := X"00000000";
		ram_buffer(7867) := X"00000000";
		ram_buffer(7868) := X"00000000";
		ram_buffer(7869) := X"00000000";
		ram_buffer(7870) := X"00000000";
		ram_buffer(7871) := X"00000000";
		ram_buffer(7872) := X"00000000";
		ram_buffer(7873) := X"00000000";
		ram_buffer(7874) := X"00000000";
		ram_buffer(7875) := X"00000000";
		ram_buffer(7876) := X"00000000";
		ram_buffer(7877) := X"00000000";
		ram_buffer(7878) := X"00000000";
		ram_buffer(7879) := X"00000000";
		ram_buffer(7880) := X"00000000";
		ram_buffer(7881) := X"00000000";
		ram_buffer(7882) := X"00000000";
		ram_buffer(7883) := X"00000000";
		ram_buffer(7884) := X"00000000";
		ram_buffer(7885) := X"00000000";
		ram_buffer(7886) := X"00000000";
		ram_buffer(7887) := X"00000000";
		ram_buffer(7888) := X"00000000";
		ram_buffer(7889) := X"00000000";
		ram_buffer(7890) := X"00000000";
		ram_buffer(7891) := X"00000000";
		ram_buffer(7892) := X"00000000";
		ram_buffer(7893) := X"00000000";
		ram_buffer(7894) := X"00000000";
		ram_buffer(7895) := X"00000000";
		ram_buffer(7896) := X"00000000";
		ram_buffer(7897) := X"00000000";
		ram_buffer(7898) := X"00000000";
		ram_buffer(7899) := X"00000000";
		ram_buffer(7900) := X"00000000";
		ram_buffer(7901) := X"00000000";
		ram_buffer(7902) := X"00000000";
		ram_buffer(7903) := X"00000000";
		ram_buffer(7904) := X"00000000";
		ram_buffer(7905) := X"00000000";
		ram_buffer(7906) := X"00000000";
		ram_buffer(7907) := X"00000000";
		ram_buffer(7908) := X"00000000";
		ram_buffer(7909) := X"00000000";
		ram_buffer(7910) := X"00000000";
		ram_buffer(7911) := X"00000000";
		ram_buffer(7912) := X"00000000";
		ram_buffer(7913) := X"00000000";
		ram_buffer(7914) := X"00000000";
		ram_buffer(7915) := X"00000000";
		ram_buffer(7916) := X"00000000";
		ram_buffer(7917) := X"00000000";
		ram_buffer(7918) := X"00000000";
		ram_buffer(7919) := X"00000000";
		ram_buffer(7920) := X"00000000";
		ram_buffer(7921) := X"00000000";
		ram_buffer(7922) := X"00000000";
		ram_buffer(7923) := X"00000000";
		ram_buffer(7924) := X"00000000";
		ram_buffer(7925) := X"00000000";
		ram_buffer(7926) := X"00000000";
		ram_buffer(7927) := X"00000000";
		ram_buffer(7928) := X"00000000";
		ram_buffer(7929) := X"00000000";
		ram_buffer(7930) := X"00000000";
		ram_buffer(7931) := X"00000000";
		ram_buffer(7932) := X"00000000";
		ram_buffer(7933) := X"00000000";
		ram_buffer(7934) := X"00000000";
		ram_buffer(7935) := X"00000000";
		ram_buffer(7936) := X"00000000";
		ram_buffer(7937) := X"00000000";
		ram_buffer(7938) := X"00000000";
		ram_buffer(7939) := X"00000000";
		ram_buffer(7940) := X"00000000";
		ram_buffer(7941) := X"00000000";
		ram_buffer(7942) := X"00000000";
		ram_buffer(7943) := X"00000000";
		ram_buffer(7944) := X"00000000";
		ram_buffer(7945) := X"00000000";
		ram_buffer(7946) := X"00000000";
		ram_buffer(7947) := X"00000000";
		ram_buffer(7948) := X"00000000";
		ram_buffer(7949) := X"00000000";
		ram_buffer(7950) := X"00000000";
		ram_buffer(7951) := X"00000000";
		ram_buffer(7952) := X"00000000";
		ram_buffer(7953) := X"00000000";
		ram_buffer(7954) := X"00000000";
		ram_buffer(7955) := X"00000000";
		ram_buffer(7956) := X"00000000";
		ram_buffer(7957) := X"00000000";
		ram_buffer(7958) := X"00000000";
		ram_buffer(7959) := X"00000000";
		ram_buffer(7960) := X"00000000";
		ram_buffer(7961) := X"00000000";
		ram_buffer(7962) := X"00000000";
		ram_buffer(7963) := X"00000000";
		ram_buffer(7964) := X"00000000";
		ram_buffer(7965) := X"00000000";
		ram_buffer(7966) := X"00000000";
		ram_buffer(7967) := X"00000000";
		ram_buffer(7968) := X"00000000";
		ram_buffer(7969) := X"00000000";
		ram_buffer(7970) := X"00000000";
		ram_buffer(7971) := X"00000000";
		ram_buffer(7972) := X"00000000";
		ram_buffer(7973) := X"00000000";
		ram_buffer(7974) := X"00000000";
		ram_buffer(7975) := X"00000000";
		ram_buffer(7976) := X"00000000";
		ram_buffer(7977) := X"00000000";
		ram_buffer(7978) := X"00000000";
		ram_buffer(7979) := X"00000000";
		ram_buffer(7980) := X"00000000";
		ram_buffer(7981) := X"00000000";
		ram_buffer(7982) := X"00000000";
		ram_buffer(7983) := X"00000000";
		ram_buffer(7984) := X"00000000";
		ram_buffer(7985) := X"00000000";
		ram_buffer(7986) := X"00000000";
		ram_buffer(7987) := X"00000000";
		ram_buffer(7988) := X"00000000";
		ram_buffer(7989) := X"00000000";
		ram_buffer(7990) := X"00000000";
		ram_buffer(7991) := X"00000000";
		ram_buffer(7992) := X"00000000";
		ram_buffer(7993) := X"00000000";
		ram_buffer(7994) := X"00000000";
		ram_buffer(7995) := X"00000000";
		ram_buffer(7996) := X"00000000";
		ram_buffer(7997) := X"00000000";
		ram_buffer(7998) := X"00000000";
		ram_buffer(7999) := X"00000000";
		ram_buffer(8000) := X"00000000";
		ram_buffer(8001) := X"00000000";
		ram_buffer(8002) := X"00000000";
		ram_buffer(8003) := X"00000000";
		ram_buffer(8004) := X"00000000";
		ram_buffer(8005) := X"00000000";
		ram_buffer(8006) := X"00000000";
		ram_buffer(8007) := X"00000000";
		ram_buffer(8008) := X"00000000";
		ram_buffer(8009) := X"00000000";
		ram_buffer(8010) := X"00000000";
		ram_buffer(8011) := X"00000000";
		ram_buffer(8012) := X"00000000";
		ram_buffer(8013) := X"00000000";
		ram_buffer(8014) := X"00000000";
		ram_buffer(8015) := X"00000000";
		ram_buffer(8016) := X"00000000";
		ram_buffer(8017) := X"00000000";
		ram_buffer(8018) := X"00000000";
		ram_buffer(8019) := X"00000000";
		ram_buffer(8020) := X"00000000";
		ram_buffer(8021) := X"00000000";
		ram_buffer(8022) := X"00000000";
		ram_buffer(8023) := X"00000000";
		ram_buffer(8024) := X"00000000";
		ram_buffer(8025) := X"00000000";
		ram_buffer(8026) := X"00000000";
		ram_buffer(8027) := X"00000000";
		ram_buffer(8028) := X"00000000";
		ram_buffer(8029) := X"00000000";
		ram_buffer(8030) := X"00000000";
		ram_buffer(8031) := X"00000000";
		ram_buffer(8032) := X"00000000";
		ram_buffer(8033) := X"00000000";
		ram_buffer(8034) := X"00000000";
		ram_buffer(8035) := X"00000000";
		ram_buffer(8036) := X"00000000";
		ram_buffer(8037) := X"00000000";
		ram_buffer(8038) := X"00000000";
		ram_buffer(8039) := X"00000000";
		ram_buffer(8040) := X"00000000";
		ram_buffer(8041) := X"00000000";
		ram_buffer(8042) := X"00000000";
		ram_buffer(8043) := X"00000000";
		ram_buffer(8044) := X"00000000";
		ram_buffer(8045) := X"00000000";
		ram_buffer(8046) := X"00000000";
		ram_buffer(8047) := X"00000000";
		ram_buffer(8048) := X"00000000";
		ram_buffer(8049) := X"00000000";
		ram_buffer(8050) := X"00000000";
		ram_buffer(8051) := X"00000000";
		ram_buffer(8052) := X"00000000";
		ram_buffer(8053) := X"00000000";
		ram_buffer(8054) := X"00000000";
		ram_buffer(8055) := X"00000000";
		ram_buffer(8056) := X"00000000";
		ram_buffer(8057) := X"00000000";
		ram_buffer(8058) := X"00000000";
		ram_buffer(8059) := X"00000000";
		ram_buffer(8060) := X"00000000";
		ram_buffer(8061) := X"00000000";
		ram_buffer(8062) := X"00000000";
		ram_buffer(8063) := X"00000000";
		ram_buffer(8064) := X"00000000";
		ram_buffer(8065) := X"00000000";
		ram_buffer(8066) := X"00000000";
		ram_buffer(8067) := X"00000000";
		ram_buffer(8068) := X"00000000";
		ram_buffer(8069) := X"00000000";
		ram_buffer(8070) := X"00000000";
		ram_buffer(8071) := X"00000000";
		ram_buffer(8072) := X"00000000";
		ram_buffer(8073) := X"00000000";
		ram_buffer(8074) := X"00000000";
		ram_buffer(8075) := X"00000000";
		ram_buffer(8076) := X"00000000";
		ram_buffer(8077) := X"00000000";
		ram_buffer(8078) := X"00000000";
		ram_buffer(8079) := X"00000000";
		ram_buffer(8080) := X"00000000";
		ram_buffer(8081) := X"00000000";
		ram_buffer(8082) := X"00000000";
		ram_buffer(8083) := X"00000000";
		ram_buffer(8084) := X"00000000";
		ram_buffer(8085) := X"00000000";
		ram_buffer(8086) := X"00000000";
		ram_buffer(8087) := X"00000000";
		ram_buffer(8088) := X"00000000";
		ram_buffer(8089) := X"00000000";
		ram_buffer(8090) := X"00000000";
		ram_buffer(8091) := X"00000000";
		ram_buffer(8092) := X"00000000";
		ram_buffer(8093) := X"00000000";
		ram_buffer(8094) := X"00000000";
		ram_buffer(8095) := X"00000000";
		ram_buffer(8096) := X"00000000";
		ram_buffer(8097) := X"00000000";
		ram_buffer(8098) := X"00000000";
		ram_buffer(8099) := X"00000000";
		ram_buffer(8100) := X"00000000";
		ram_buffer(8101) := X"00000000";
		ram_buffer(8102) := X"00000000";
		ram_buffer(8103) := X"00000000";
		ram_buffer(8104) := X"00000000";
		ram_buffer(8105) := X"00000000";
		ram_buffer(8106) := X"00000000";
		ram_buffer(8107) := X"00000000";
		ram_buffer(8108) := X"00000000";
		ram_buffer(8109) := X"00000000";
		ram_buffer(8110) := X"00000000";
		ram_buffer(8111) := X"00000000";
		ram_buffer(8112) := X"00000000";
		ram_buffer(8113) := X"00000000";
		ram_buffer(8114) := X"00000000";
		ram_buffer(8115) := X"00000000";
		ram_buffer(8116) := X"00000000";
		ram_buffer(8117) := X"00000000";
		ram_buffer(8118) := X"00000000";
		ram_buffer(8119) := X"00000000";
		ram_buffer(8120) := X"00000000";
		ram_buffer(8121) := X"00000000";
		ram_buffer(8122) := X"00000000";
		ram_buffer(8123) := X"00000000";
		ram_buffer(8124) := X"00000000";
		ram_buffer(8125) := X"00000000";
		ram_buffer(8126) := X"00000000";
		ram_buffer(8127) := X"00000000";
		ram_buffer(8128) := X"00000000";
		ram_buffer(8129) := X"00000000";
		ram_buffer(8130) := X"00000000";
		ram_buffer(8131) := X"00000000";
		ram_buffer(8132) := X"00000000";
		ram_buffer(8133) := X"00000000";
		ram_buffer(8134) := X"00000000";
		ram_buffer(8135) := X"00000000";
		ram_buffer(8136) := X"00000000";
		ram_buffer(8137) := X"00000000";
		ram_buffer(8138) := X"00000000";
		ram_buffer(8139) := X"00000000";
		ram_buffer(8140) := X"00000000";
		ram_buffer(8141) := X"00000000";
		ram_buffer(8142) := X"00000000";
		ram_buffer(8143) := X"00000000";
		ram_buffer(8144) := X"00000000";
		ram_buffer(8145) := X"00000000";
		ram_buffer(8146) := X"00000000";
		ram_buffer(8147) := X"00000000";
		ram_buffer(8148) := X"00000000";
		ram_buffer(8149) := X"00000000";
		ram_buffer(8150) := X"00000000";
		ram_buffer(8151) := X"00000000";
		ram_buffer(8152) := X"00000000";
		ram_buffer(8153) := X"00000000";
		ram_buffer(8154) := X"00000000";
		ram_buffer(8155) := X"00000000";
		ram_buffer(8156) := X"00000000";
		ram_buffer(8157) := X"00000000";
		ram_buffer(8158) := X"00000000";
		ram_buffer(8159) := X"00000000";
		ram_buffer(8160) := X"00000000";
		ram_buffer(8161) := X"00000000";
		ram_buffer(8162) := X"00000000";
		ram_buffer(8163) := X"00000000";
		ram_buffer(8164) := X"00000000";
		ram_buffer(8165) := X"00000000";
		ram_buffer(8166) := X"00000000";
		ram_buffer(8167) := X"00000000";
		ram_buffer(8168) := X"00000000";
		ram_buffer(8169) := X"00000000";
		ram_buffer(8170) := X"00000000";
		ram_buffer(8171) := X"00000000";
		ram_buffer(8172) := X"00000000";
		ram_buffer(8173) := X"00000000";
		ram_buffer(8174) := X"00000000";
		ram_buffer(8175) := X"00000000";
		ram_buffer(8176) := X"00000000";
		ram_buffer(8177) := X"00000000";
		ram_buffer(8178) := X"00000000";
		ram_buffer(8179) := X"00000000";
		ram_buffer(8180) := X"00000000";
		ram_buffer(8181) := X"00000000";
		ram_buffer(8182) := X"00000000";
		ram_buffer(8183) := X"00000000";
		ram_buffer(8184) := X"00000000";
		ram_buffer(8185) := X"00000000";
		ram_buffer(8186) := X"00000000";
		ram_buffer(8187) := X"00000000";
		ram_buffer(8188) := X"00000000";
		ram_buffer(8189) := X"00000000";
		ram_buffer(8190) := X"00000000";
		ram_buffer(8191) := X"00000000";
		return ram_buffer;
	end;
end;
