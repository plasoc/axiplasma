library ieee;
use ieee.std_logic_1164.all;

package bram_pack is

	constant cpu_width : integer := 32;
	constant ram_size : integer := 16384;
	subtype word_type is std_logic_vector(cpu_width-1 downto 0);
	type ram_type is array(0 to ram_size-1) of word_type;
	function load_hex return ram_type;

end package;

package body bram_pack is

	function load_hex return ram_type is
		variable ram_buffer : ram_type;
	begin
		ram_buffer(0) := X"3C1C0001";
		ram_buffer(1) := X"279C83F0";
		ram_buffer(2) := X"3C050000";
		ram_buffer(3) := X"24A503FC";
		ram_buffer(4) := X"3C040000";
		ram_buffer(5) := X"24840654";
		ram_buffer(6) := X"3C1D0000";
		ram_buffer(7) := X"27BD05F8";
		ram_buffer(8) := X"ACA00000";
		ram_buffer(9) := X"00A4182A";
		ram_buffer(10) := X"1460FFFD";
		ram_buffer(11) := X"24A50004";
		ram_buffer(12) := X"0C00007C";
		ram_buffer(13) := X"00000000";
		ram_buffer(14) := X"0800000E";
		ram_buffer(15) := X"23BDFF98";
		ram_buffer(16) := X"AFA10010";
		ram_buffer(17) := X"AFA20014";
		ram_buffer(18) := X"AFA30018";
		ram_buffer(19) := X"AFA4001C";
		ram_buffer(20) := X"AFA50020";
		ram_buffer(21) := X"AFA60024";
		ram_buffer(22) := X"AFA70028";
		ram_buffer(23) := X"AFA8002C";
		ram_buffer(24) := X"AFA90030";
		ram_buffer(25) := X"AFAA0034";
		ram_buffer(26) := X"AFAB0038";
		ram_buffer(27) := X"AFAC003C";
		ram_buffer(28) := X"AFAD0040";
		ram_buffer(29) := X"AFAE0044";
		ram_buffer(30) := X"AFAF0048";
		ram_buffer(31) := X"AFB8004C";
		ram_buffer(32) := X"AFB90050";
		ram_buffer(33) := X"AFBF0054";
		ram_buffer(34) := X"401A7000";
		ram_buffer(35) := X"235AFFFC";
		ram_buffer(36) := X"AFBA0058";
		ram_buffer(37) := X"0000D810";
		ram_buffer(38) := X"AFBB005C";
		ram_buffer(39) := X"0000D812";
		ram_buffer(40) := X"AFBB0060";
		ram_buffer(41) := X"0C0000CC";
		ram_buffer(42) := X"23A50000";
		ram_buffer(43) := X"8FA10010";
		ram_buffer(44) := X"8FA20014";
		ram_buffer(45) := X"8FA30018";
		ram_buffer(46) := X"8FA4001C";
		ram_buffer(47) := X"8FA50020";
		ram_buffer(48) := X"8FA60024";
		ram_buffer(49) := X"8FA70028";
		ram_buffer(50) := X"8FA8002C";
		ram_buffer(51) := X"8FA90030";
		ram_buffer(52) := X"8FAA0034";
		ram_buffer(53) := X"8FAB0038";
		ram_buffer(54) := X"8FAC003C";
		ram_buffer(55) := X"8FAD0040";
		ram_buffer(56) := X"8FAE0044";
		ram_buffer(57) := X"8FAF0048";
		ram_buffer(58) := X"8FB8004C";
		ram_buffer(59) := X"8FB90050";
		ram_buffer(60) := X"8FBF0054";
		ram_buffer(61) := X"8FBA0058";
		ram_buffer(62) := X"8FBB005C";
		ram_buffer(63) := X"03600011";
		ram_buffer(64) := X"8FBB0060";
		ram_buffer(65) := X"03600013";
		ram_buffer(66) := X"23BD0068";
		ram_buffer(67) := X"341B0001";
		ram_buffer(68) := X"03400008";
		ram_buffer(69) := X"409B6000";
		ram_buffer(70) := X"40026000";
		ram_buffer(71) := X"03E00008";
		ram_buffer(72) := X"40846000";
		ram_buffer(73) := X"3C050000";
		ram_buffer(74) := X"24A50150";
		ram_buffer(75) := X"8CA60000";
		ram_buffer(76) := X"AC06003C";
		ram_buffer(77) := X"8CA60004";
		ram_buffer(78) := X"AC060040";
		ram_buffer(79) := X"8CA60008";
		ram_buffer(80) := X"AC060044";
		ram_buffer(81) := X"8CA6000C";
		ram_buffer(82) := X"03E00008";
		ram_buffer(83) := X"AC060048";
		ram_buffer(84) := X"3C1A1000";
		ram_buffer(85) := X"375A003C";
		ram_buffer(86) := X"03400008";
		ram_buffer(87) := X"00000000";
		ram_buffer(88) := X"AC900000";
		ram_buffer(89) := X"AC910004";
		ram_buffer(90) := X"AC920008";
		ram_buffer(91) := X"AC93000C";
		ram_buffer(92) := X"AC940010";
		ram_buffer(93) := X"AC950014";
		ram_buffer(94) := X"AC960018";
		ram_buffer(95) := X"AC97001C";
		ram_buffer(96) := X"AC9E0020";
		ram_buffer(97) := X"AC9C0024";
		ram_buffer(98) := X"AC9D0028";
		ram_buffer(99) := X"AC9F002C";
		ram_buffer(100) := X"03E00008";
		ram_buffer(101) := X"34020000";
		ram_buffer(102) := X"8C900000";
		ram_buffer(103) := X"8C910004";
		ram_buffer(104) := X"8C920008";
		ram_buffer(105) := X"8C93000C";
		ram_buffer(106) := X"8C940010";
		ram_buffer(107) := X"8C950014";
		ram_buffer(108) := X"8C960018";
		ram_buffer(109) := X"8C97001C";
		ram_buffer(110) := X"8C9E0020";
		ram_buffer(111) := X"8C9C0024";
		ram_buffer(112) := X"8C9D0028";
		ram_buffer(113) := X"8C9F002C";
		ram_buffer(114) := X"03E00008";
		ram_buffer(115) := X"34A20000";
		ram_buffer(116) := X"00850019";
		ram_buffer(117) := X"00001012";
		ram_buffer(118) := X"00002010";
		ram_buffer(119) := X"03E00008";
		ram_buffer(120) := X"ACC40000";
		ram_buffer(121) := X"0000000C";
		ram_buffer(122) := X"03E00008";
		ram_buffer(123) := X"00000000";
		ram_buffer(124) := X"27BDFFE8";
		ram_buffer(125) := X"3C0344A0";
		ram_buffer(126) := X"AFB00010";
		ram_buffer(127) := X"3C100000";
		ram_buffer(128) := X"AE030610";
		ram_buffer(129) := X"3C0344A2";
		ram_buffer(130) := X"AF838014";
		ram_buffer(131) := X"3C03017D";
		ram_buffer(132) := X"3C0444A1";
		ram_buffer(133) := X"24637840";
		ram_buffer(134) := X"AFBF0014";
		ram_buffer(135) := X"AF848010";
		ram_buffer(136) := X"AC830004";
		ram_buffer(137) := X"3C030000";
		ram_buffer(138) := X"26020610";
		ram_buffer(139) := X"24630304";
		ram_buffer(140) := X"AC43000C";
		ram_buffer(141) := X"3C030000";
		ram_buffer(142) := X"246302DC";
		ram_buffer(143) := X"24040001";
		ram_buffer(144) := X"AC430004";
		ram_buffer(145) := X"AC400014";
		ram_buffer(146) := X"AC40001C";
		ram_buffer(147) := X"AC400024";
		ram_buffer(148) := X"AC40002C";
		ram_buffer(149) := X"AC400034";
		ram_buffer(150) := X"AC40003C";
		ram_buffer(151) := X"AC400010";
		ram_buffer(152) := X"0C000046";
		ram_buffer(153) := X"AC400008";
		ram_buffer(154) := X"8E020610";
		ram_buffer(155) := X"240300FF";
		ram_buffer(156) := X"AC430000";
		ram_buffer(157) := X"8F828010";
		ram_buffer(158) := X"24030003";
		ram_buffer(159) := X"AC430000";
		ram_buffer(160) := X"8F828014";
		ram_buffer(161) := X"24030001";
		ram_buffer(162) := X"AC430000";
		ram_buffer(163) := X"240400FF";
		ram_buffer(164) := X"8F828008";
		ram_buffer(165) := X"00000000";
		ram_buffer(166) := X"1040FFFD";
		ram_buffer(167) := X"00000000";
		ram_buffer(168) := X"8E020610";
		ram_buffer(169) := X"00000000";
		ram_buffer(170) := X"AC400000";
		ram_buffer(171) := X"AF808008";
		ram_buffer(172) := X"8F828018";
		ram_buffer(173) := X"8F83800C";
		ram_buffer(174) := X"00000000";
		ram_buffer(175) := X"00430018";
		ram_buffer(176) := X"8F838014";
		ram_buffer(177) := X"00001012";
		ram_buffer(178) := X"AC620008";
		ram_buffer(179) := X"8E020610";
		ram_buffer(180) := X"00000000";
		ram_buffer(181) := X"1000FFEE";
		ram_buffer(182) := X"AC440000";
		ram_buffer(183) := X"8F82800C";
		ram_buffer(184) := X"00000000";
		ram_buffer(185) := X"2C420001";
		ram_buffer(186) := X"AF82800C";
		ram_buffer(187) := X"24020001";
		ram_buffer(188) := X"AF828008";
		ram_buffer(189) := X"8F828010";
		ram_buffer(190) := X"24030007";
		ram_buffer(191) := X"03E00008";
		ram_buffer(192) := X"AC430000";
		ram_buffer(193) := X"8F838014";
		ram_buffer(194) := X"24020001";
		ram_buffer(195) := X"8C630004";
		ram_buffer(196) := X"00000000";
		ram_buffer(197) := X"AF838018";
		ram_buffer(198) := X"AF82800C";
		ram_buffer(199) := X"AF828008";
		ram_buffer(200) := X"8F828014";
		ram_buffer(201) := X"24030003";
		ram_buffer(202) := X"03E00008";
		ram_buffer(203) := X"AC430000";
		ram_buffer(204) := X"27BDFFE0";
		ram_buffer(205) := X"AFB10018";
		ram_buffer(206) := X"3C110000";
		ram_buffer(207) := X"8E220610";
		ram_buffer(208) := X"AFBF001C";
		ram_buffer(209) := X"8C420004";
		ram_buffer(210) := X"00000000";
		ram_buffer(211) := X"2C430008";
		ram_buffer(212) := X"10600010";
		ram_buffer(213) := X"AFB00014";
		ram_buffer(214) := X"3C100000";
		ram_buffer(215) := X"26100614";
		ram_buffer(216) := X"000210C0";
		ram_buffer(217) := X"02021021";
		ram_buffer(218) := X"8C430000";
		ram_buffer(219) := X"8C440004";
		ram_buffer(220) := X"0060F809";
		ram_buffer(221) := X"00000000";
		ram_buffer(222) := X"8E220610";
		ram_buffer(223) := X"00000000";
		ram_buffer(224) := X"8C420004";
		ram_buffer(225) := X"00000000";
		ram_buffer(226) := X"2C430008";
		ram_buffer(227) := X"1460FFF4";
		ram_buffer(228) := X"00000000";
		ram_buffer(229) := X"8FBF001C";
		ram_buffer(230) := X"8FB10018";
		ram_buffer(231) := X"8FB00014";
		ram_buffer(232) := X"03E00008";
		ram_buffer(233) := X"27BD0020";
		ram_buffer(234) := X"10C00011";
		ram_buffer(235) := X"00C51821";
		ram_buffer(236) := X"2406FFE0";
		ram_buffer(237) := X"00661024";
		ram_buffer(238) := X"0043182B";
		ram_buffer(239) := X"00031940";
		ram_buffer(240) := X"24420020";
		ram_buffer(241) := X"00A62824";
		ram_buffer(242) := X"00431821";
		ram_buffer(243) := X"10A30008";
		ram_buffer(244) := X"3C021000";
		ram_buffer(245) := X"00822021";
		ram_buffer(246) := X"00A61024";
		ram_buffer(247) := X"AC820000";
		ram_buffer(248) := X"AC400000";
		ram_buffer(249) := X"24A50020";
		ram_buffer(250) := X"14A3FFFC";
		ram_buffer(251) := X"00A61024";
		ram_buffer(252) := X"03E00008";
		ram_buffer(253) := X"00000000";
		ram_buffer(254) := X"00000001";
		ram_buffer(255) := X"00000000";
		ram_buffer(256) := X"00000000";
		ram_buffer(257) := X"00000000";
		ram_buffer(258) := X"00000000";
		ram_buffer(259) := X"00000000";
		ram_buffer(260) := X"00000000";
		ram_buffer(261) := X"00000000";
		ram_buffer(262) := X"00000000";
		ram_buffer(263) := X"00000000";
		ram_buffer(264) := X"00000000";
		ram_buffer(265) := X"00000000";
		ram_buffer(266) := X"00000000";
		ram_buffer(267) := X"00000000";
		ram_buffer(268) := X"00000000";
		ram_buffer(269) := X"00000000";
		ram_buffer(270) := X"00000000";
		ram_buffer(271) := X"00000000";
		ram_buffer(272) := X"00000000";
		ram_buffer(273) := X"00000000";
		ram_buffer(274) := X"00000000";
		ram_buffer(275) := X"00000000";
		ram_buffer(276) := X"00000000";
		ram_buffer(277) := X"00000000";
		ram_buffer(278) := X"00000000";
		ram_buffer(279) := X"00000000";
		ram_buffer(280) := X"00000000";
		ram_buffer(281) := X"00000000";
		ram_buffer(282) := X"00000000";
		ram_buffer(283) := X"00000000";
		ram_buffer(284) := X"00000000";
		ram_buffer(285) := X"00000000";
		ram_buffer(286) := X"00000000";
		ram_buffer(287) := X"00000000";
		ram_buffer(288) := X"00000000";
		ram_buffer(289) := X"00000000";
		ram_buffer(290) := X"00000000";
		ram_buffer(291) := X"00000000";
		ram_buffer(292) := X"00000000";
		ram_buffer(293) := X"00000000";
		ram_buffer(294) := X"00000000";
		ram_buffer(295) := X"00000000";
		ram_buffer(296) := X"00000000";
		ram_buffer(297) := X"00000000";
		ram_buffer(298) := X"00000000";
		ram_buffer(299) := X"00000000";
		ram_buffer(300) := X"00000000";
		ram_buffer(301) := X"00000000";
		ram_buffer(302) := X"00000000";
		ram_buffer(303) := X"00000000";
		ram_buffer(304) := X"00000000";
		ram_buffer(305) := X"00000000";
		ram_buffer(306) := X"00000000";
		ram_buffer(307) := X"00000000";
		ram_buffer(308) := X"00000000";
		ram_buffer(309) := X"00000000";
		ram_buffer(310) := X"00000000";
		ram_buffer(311) := X"00000000";
		ram_buffer(312) := X"00000000";
		ram_buffer(313) := X"00000000";
		ram_buffer(314) := X"00000000";
		ram_buffer(315) := X"00000000";
		ram_buffer(316) := X"00000000";
		ram_buffer(317) := X"00000000";
		ram_buffer(318) := X"00000000";
		ram_buffer(319) := X"00000000";
		ram_buffer(320) := X"00000000";
		ram_buffer(321) := X"00000000";
		ram_buffer(322) := X"00000000";
		ram_buffer(323) := X"00000000";
		ram_buffer(324) := X"00000000";
		ram_buffer(325) := X"00000000";
		ram_buffer(326) := X"00000000";
		ram_buffer(327) := X"00000000";
		ram_buffer(328) := X"00000000";
		ram_buffer(329) := X"00000000";
		ram_buffer(330) := X"00000000";
		ram_buffer(331) := X"00000000";
		ram_buffer(332) := X"00000000";
		ram_buffer(333) := X"00000000";
		ram_buffer(334) := X"00000000";
		ram_buffer(335) := X"00000000";
		ram_buffer(336) := X"00000000";
		ram_buffer(337) := X"00000000";
		ram_buffer(338) := X"00000000";
		ram_buffer(339) := X"00000000";
		ram_buffer(340) := X"00000000";
		ram_buffer(341) := X"00000000";
		ram_buffer(342) := X"00000000";
		ram_buffer(343) := X"00000000";
		ram_buffer(344) := X"00000000";
		ram_buffer(345) := X"00000000";
		ram_buffer(346) := X"00000000";
		ram_buffer(347) := X"00000000";
		ram_buffer(348) := X"00000000";
		ram_buffer(349) := X"00000000";
		ram_buffer(350) := X"00000000";
		ram_buffer(351) := X"00000000";
		ram_buffer(352) := X"00000000";
		ram_buffer(353) := X"00000000";
		ram_buffer(354) := X"00000000";
		ram_buffer(355) := X"00000000";
		ram_buffer(356) := X"00000000";
		ram_buffer(357) := X"00000000";
		ram_buffer(358) := X"00000000";
		ram_buffer(359) := X"00000000";
		ram_buffer(360) := X"00000000";
		ram_buffer(361) := X"00000000";
		ram_buffer(362) := X"00000000";
		ram_buffer(363) := X"00000000";
		ram_buffer(364) := X"00000000";
		ram_buffer(365) := X"00000000";
		ram_buffer(366) := X"00000000";
		ram_buffer(367) := X"00000000";
		ram_buffer(368) := X"00000000";
		ram_buffer(369) := X"00000000";
		ram_buffer(370) := X"00000000";
		ram_buffer(371) := X"00000000";
		ram_buffer(372) := X"00000000";
		ram_buffer(373) := X"00000000";
		ram_buffer(374) := X"00000000";
		ram_buffer(375) := X"00000000";
		ram_buffer(376) := X"00000000";
		ram_buffer(377) := X"00000000";
		ram_buffer(378) := X"00000000";
		ram_buffer(379) := X"00000000";
		ram_buffer(380) := X"00000000";
		ram_buffer(381) := X"00000000";
		ram_buffer(382) := X"00000000";
		ram_buffer(383) := X"00000000";
		ram_buffer(384) := X"00000000";
		ram_buffer(385) := X"00000000";
		ram_buffer(386) := X"00000000";
		ram_buffer(387) := X"00000000";
		ram_buffer(388) := X"00000000";
		ram_buffer(389) := X"00000000";
		ram_buffer(390) := X"00000000";
		ram_buffer(391) := X"00000000";
		ram_buffer(392) := X"00000000";
		ram_buffer(393) := X"00000000";
		ram_buffer(394) := X"00000000";
		ram_buffer(395) := X"00000000";
		ram_buffer(396) := X"00000000";
		ram_buffer(397) := X"00000000";
		ram_buffer(398) := X"00000000";
		ram_buffer(399) := X"00000000";
		ram_buffer(400) := X"00000000";
		ram_buffer(401) := X"00000000";
		ram_buffer(402) := X"00000000";
		ram_buffer(403) := X"00000000";
		ram_buffer(404) := X"00000000";
		ram_buffer(405) := X"00000000";
		ram_buffer(406) := X"00000000";
		ram_buffer(407) := X"00000000";
		ram_buffer(408) := X"00000000";
		ram_buffer(409) := X"00000000";
		ram_buffer(410) := X"00000000";
		ram_buffer(411) := X"00000000";
		ram_buffer(412) := X"00000000";
		ram_buffer(413) := X"00000000";
		ram_buffer(414) := X"00000000";
		ram_buffer(415) := X"00000000";
		ram_buffer(416) := X"00000000";
		ram_buffer(417) := X"00000000";
		ram_buffer(418) := X"00000000";
		ram_buffer(419) := X"00000000";
		ram_buffer(420) := X"00000000";
		ram_buffer(421) := X"00000000";
		ram_buffer(422) := X"00000000";
		ram_buffer(423) := X"00000000";
		ram_buffer(424) := X"00000000";
		ram_buffer(425) := X"00000000";
		ram_buffer(426) := X"00000000";
		ram_buffer(427) := X"00000000";
		ram_buffer(428) := X"00000000";
		ram_buffer(429) := X"00000000";
		ram_buffer(430) := X"00000000";
		ram_buffer(431) := X"00000000";
		ram_buffer(432) := X"00000000";
		ram_buffer(433) := X"00000000";
		ram_buffer(434) := X"00000000";
		ram_buffer(435) := X"00000000";
		ram_buffer(436) := X"00000000";
		ram_buffer(437) := X"00000000";
		ram_buffer(438) := X"00000000";
		ram_buffer(439) := X"00000000";
		ram_buffer(440) := X"00000000";
		ram_buffer(441) := X"00000000";
		ram_buffer(442) := X"00000000";
		ram_buffer(443) := X"00000000";
		ram_buffer(444) := X"00000000";
		ram_buffer(445) := X"00000000";
		ram_buffer(446) := X"00000000";
		ram_buffer(447) := X"00000000";
		ram_buffer(448) := X"00000000";
		ram_buffer(449) := X"00000000";
		ram_buffer(450) := X"00000000";
		ram_buffer(451) := X"00000000";
		ram_buffer(452) := X"00000000";
		ram_buffer(453) := X"00000000";
		ram_buffer(454) := X"00000000";
		ram_buffer(455) := X"00000000";
		ram_buffer(456) := X"00000000";
		ram_buffer(457) := X"00000000";
		ram_buffer(458) := X"00000000";
		ram_buffer(459) := X"00000000";
		ram_buffer(460) := X"00000000";
		ram_buffer(461) := X"00000000";
		ram_buffer(462) := X"00000000";
		ram_buffer(463) := X"00000000";
		ram_buffer(464) := X"00000000";
		ram_buffer(465) := X"00000000";
		ram_buffer(466) := X"00000000";
		ram_buffer(467) := X"00000000";
		ram_buffer(468) := X"00000000";
		ram_buffer(469) := X"00000000";
		ram_buffer(470) := X"00000000";
		ram_buffer(471) := X"00000000";
		ram_buffer(472) := X"00000000";
		ram_buffer(473) := X"00000000";
		ram_buffer(474) := X"00000000";
		ram_buffer(475) := X"00000000";
		ram_buffer(476) := X"00000000";
		ram_buffer(477) := X"00000000";
		ram_buffer(478) := X"00000000";
		ram_buffer(479) := X"00000000";
		ram_buffer(480) := X"00000000";
		ram_buffer(481) := X"00000000";
		ram_buffer(482) := X"00000000";
		ram_buffer(483) := X"00000000";
		ram_buffer(484) := X"00000000";
		ram_buffer(485) := X"00000000";
		ram_buffer(486) := X"00000000";
		ram_buffer(487) := X"00000000";
		ram_buffer(488) := X"00000000";
		ram_buffer(489) := X"00000000";
		ram_buffer(490) := X"00000000";
		ram_buffer(491) := X"00000000";
		ram_buffer(492) := X"00000000";
		ram_buffer(493) := X"00000000";
		ram_buffer(494) := X"00000000";
		ram_buffer(495) := X"00000000";
		ram_buffer(496) := X"00000000";
		ram_buffer(497) := X"00000000";
		ram_buffer(498) := X"00000000";
		ram_buffer(499) := X"00000000";
		ram_buffer(500) := X"00000000";
		ram_buffer(501) := X"00000000";
		ram_buffer(502) := X"00000000";
		ram_buffer(503) := X"00000000";
		ram_buffer(504) := X"00000000";
		ram_buffer(505) := X"00000000";
		ram_buffer(506) := X"00000000";
		ram_buffer(507) := X"00000000";
		ram_buffer(508) := X"00000000";
		ram_buffer(509) := X"00000000";
		ram_buffer(510) := X"00000000";
		ram_buffer(511) := X"00000000";
		ram_buffer(512) := X"00000000";
		ram_buffer(513) := X"00000000";
		ram_buffer(514) := X"00000000";
		ram_buffer(515) := X"00000000";
		ram_buffer(516) := X"00000000";
		ram_buffer(517) := X"00000000";
		ram_buffer(518) := X"00000000";
		ram_buffer(519) := X"00000000";
		ram_buffer(520) := X"00000000";
		ram_buffer(521) := X"00000000";
		ram_buffer(522) := X"00000000";
		ram_buffer(523) := X"00000000";
		ram_buffer(524) := X"00000000";
		ram_buffer(525) := X"00000000";
		ram_buffer(526) := X"00000000";
		ram_buffer(527) := X"00000000";
		ram_buffer(528) := X"00000000";
		ram_buffer(529) := X"00000000";
		ram_buffer(530) := X"00000000";
		ram_buffer(531) := X"00000000";
		ram_buffer(532) := X"00000000";
		ram_buffer(533) := X"00000000";
		ram_buffer(534) := X"00000000";
		ram_buffer(535) := X"00000000";
		ram_buffer(536) := X"00000000";
		ram_buffer(537) := X"00000000";
		ram_buffer(538) := X"00000000";
		ram_buffer(539) := X"00000000";
		ram_buffer(540) := X"00000000";
		ram_buffer(541) := X"00000000";
		ram_buffer(542) := X"00000000";
		ram_buffer(543) := X"00000000";
		ram_buffer(544) := X"00000000";
		ram_buffer(545) := X"00000000";
		ram_buffer(546) := X"00000000";
		ram_buffer(547) := X"00000000";
		ram_buffer(548) := X"00000000";
		ram_buffer(549) := X"00000000";
		ram_buffer(550) := X"00000000";
		ram_buffer(551) := X"00000000";
		ram_buffer(552) := X"00000000";
		ram_buffer(553) := X"00000000";
		ram_buffer(554) := X"00000000";
		ram_buffer(555) := X"00000000";
		ram_buffer(556) := X"00000000";
		ram_buffer(557) := X"00000000";
		ram_buffer(558) := X"00000000";
		ram_buffer(559) := X"00000000";
		ram_buffer(560) := X"00000000";
		ram_buffer(561) := X"00000000";
		ram_buffer(562) := X"00000000";
		ram_buffer(563) := X"00000000";
		ram_buffer(564) := X"00000000";
		ram_buffer(565) := X"00000000";
		ram_buffer(566) := X"00000000";
		ram_buffer(567) := X"00000000";
		ram_buffer(568) := X"00000000";
		ram_buffer(569) := X"00000000";
		ram_buffer(570) := X"00000000";
		ram_buffer(571) := X"00000000";
		ram_buffer(572) := X"00000000";
		ram_buffer(573) := X"00000000";
		ram_buffer(574) := X"00000000";
		ram_buffer(575) := X"00000000";
		ram_buffer(576) := X"00000000";
		ram_buffer(577) := X"00000000";
		ram_buffer(578) := X"00000000";
		ram_buffer(579) := X"00000000";
		ram_buffer(580) := X"00000000";
		ram_buffer(581) := X"00000000";
		ram_buffer(582) := X"00000000";
		ram_buffer(583) := X"00000000";
		ram_buffer(584) := X"00000000";
		ram_buffer(585) := X"00000000";
		ram_buffer(586) := X"00000000";
		ram_buffer(587) := X"00000000";
		ram_buffer(588) := X"00000000";
		ram_buffer(589) := X"00000000";
		ram_buffer(590) := X"00000000";
		ram_buffer(591) := X"00000000";
		ram_buffer(592) := X"00000000";
		ram_buffer(593) := X"00000000";
		ram_buffer(594) := X"00000000";
		ram_buffer(595) := X"00000000";
		ram_buffer(596) := X"00000000";
		ram_buffer(597) := X"00000000";
		ram_buffer(598) := X"00000000";
		ram_buffer(599) := X"00000000";
		ram_buffer(600) := X"00000000";
		ram_buffer(601) := X"00000000";
		ram_buffer(602) := X"00000000";
		ram_buffer(603) := X"00000000";
		ram_buffer(604) := X"00000000";
		ram_buffer(605) := X"00000000";
		ram_buffer(606) := X"00000000";
		ram_buffer(607) := X"00000000";
		ram_buffer(608) := X"00000000";
		ram_buffer(609) := X"00000000";
		ram_buffer(610) := X"00000000";
		ram_buffer(611) := X"00000000";
		ram_buffer(612) := X"00000000";
		ram_buffer(613) := X"00000000";
		ram_buffer(614) := X"00000000";
		ram_buffer(615) := X"00000000";
		ram_buffer(616) := X"00000000";
		ram_buffer(617) := X"00000000";
		ram_buffer(618) := X"00000000";
		ram_buffer(619) := X"00000000";
		ram_buffer(620) := X"00000000";
		ram_buffer(621) := X"00000000";
		ram_buffer(622) := X"00000000";
		ram_buffer(623) := X"00000000";
		ram_buffer(624) := X"00000000";
		ram_buffer(625) := X"00000000";
		ram_buffer(626) := X"00000000";
		ram_buffer(627) := X"00000000";
		ram_buffer(628) := X"00000000";
		ram_buffer(629) := X"00000000";
		ram_buffer(630) := X"00000000";
		ram_buffer(631) := X"00000000";
		ram_buffer(632) := X"00000000";
		ram_buffer(633) := X"00000000";
		ram_buffer(634) := X"00000000";
		ram_buffer(635) := X"00000000";
		ram_buffer(636) := X"00000000";
		ram_buffer(637) := X"00000000";
		ram_buffer(638) := X"00000000";
		ram_buffer(639) := X"00000000";
		ram_buffer(640) := X"00000000";
		ram_buffer(641) := X"00000000";
		ram_buffer(642) := X"00000000";
		ram_buffer(643) := X"00000000";
		ram_buffer(644) := X"00000000";
		ram_buffer(645) := X"00000000";
		ram_buffer(646) := X"00000000";
		ram_buffer(647) := X"00000000";
		ram_buffer(648) := X"00000000";
		ram_buffer(649) := X"00000000";
		ram_buffer(650) := X"00000000";
		ram_buffer(651) := X"00000000";
		ram_buffer(652) := X"00000000";
		ram_buffer(653) := X"00000000";
		ram_buffer(654) := X"00000000";
		ram_buffer(655) := X"00000000";
		ram_buffer(656) := X"00000000";
		ram_buffer(657) := X"00000000";
		ram_buffer(658) := X"00000000";
		ram_buffer(659) := X"00000000";
		ram_buffer(660) := X"00000000";
		ram_buffer(661) := X"00000000";
		ram_buffer(662) := X"00000000";
		ram_buffer(663) := X"00000000";
		ram_buffer(664) := X"00000000";
		ram_buffer(665) := X"00000000";
		ram_buffer(666) := X"00000000";
		ram_buffer(667) := X"00000000";
		ram_buffer(668) := X"00000000";
		ram_buffer(669) := X"00000000";
		ram_buffer(670) := X"00000000";
		ram_buffer(671) := X"00000000";
		ram_buffer(672) := X"00000000";
		ram_buffer(673) := X"00000000";
		ram_buffer(674) := X"00000000";
		ram_buffer(675) := X"00000000";
		ram_buffer(676) := X"00000000";
		ram_buffer(677) := X"00000000";
		ram_buffer(678) := X"00000000";
		ram_buffer(679) := X"00000000";
		ram_buffer(680) := X"00000000";
		ram_buffer(681) := X"00000000";
		ram_buffer(682) := X"00000000";
		ram_buffer(683) := X"00000000";
		ram_buffer(684) := X"00000000";
		ram_buffer(685) := X"00000000";
		ram_buffer(686) := X"00000000";
		ram_buffer(687) := X"00000000";
		ram_buffer(688) := X"00000000";
		ram_buffer(689) := X"00000000";
		ram_buffer(690) := X"00000000";
		ram_buffer(691) := X"00000000";
		ram_buffer(692) := X"00000000";
		ram_buffer(693) := X"00000000";
		ram_buffer(694) := X"00000000";
		ram_buffer(695) := X"00000000";
		ram_buffer(696) := X"00000000";
		ram_buffer(697) := X"00000000";
		ram_buffer(698) := X"00000000";
		ram_buffer(699) := X"00000000";
		ram_buffer(700) := X"00000000";
		ram_buffer(701) := X"00000000";
		ram_buffer(702) := X"00000000";
		ram_buffer(703) := X"00000000";
		ram_buffer(704) := X"00000000";
		ram_buffer(705) := X"00000000";
		ram_buffer(706) := X"00000000";
		ram_buffer(707) := X"00000000";
		ram_buffer(708) := X"00000000";
		ram_buffer(709) := X"00000000";
		ram_buffer(710) := X"00000000";
		ram_buffer(711) := X"00000000";
		ram_buffer(712) := X"00000000";
		ram_buffer(713) := X"00000000";
		ram_buffer(714) := X"00000000";
		ram_buffer(715) := X"00000000";
		ram_buffer(716) := X"00000000";
		ram_buffer(717) := X"00000000";
		ram_buffer(718) := X"00000000";
		ram_buffer(719) := X"00000000";
		ram_buffer(720) := X"00000000";
		ram_buffer(721) := X"00000000";
		ram_buffer(722) := X"00000000";
		ram_buffer(723) := X"00000000";
		ram_buffer(724) := X"00000000";
		ram_buffer(725) := X"00000000";
		ram_buffer(726) := X"00000000";
		ram_buffer(727) := X"00000000";
		ram_buffer(728) := X"00000000";
		ram_buffer(729) := X"00000000";
		ram_buffer(730) := X"00000000";
		ram_buffer(731) := X"00000000";
		ram_buffer(732) := X"00000000";
		ram_buffer(733) := X"00000000";
		ram_buffer(734) := X"00000000";
		ram_buffer(735) := X"00000000";
		ram_buffer(736) := X"00000000";
		ram_buffer(737) := X"00000000";
		ram_buffer(738) := X"00000000";
		ram_buffer(739) := X"00000000";
		ram_buffer(740) := X"00000000";
		ram_buffer(741) := X"00000000";
		ram_buffer(742) := X"00000000";
		ram_buffer(743) := X"00000000";
		ram_buffer(744) := X"00000000";
		ram_buffer(745) := X"00000000";
		ram_buffer(746) := X"00000000";
		ram_buffer(747) := X"00000000";
		ram_buffer(748) := X"00000000";
		ram_buffer(749) := X"00000000";
		ram_buffer(750) := X"00000000";
		ram_buffer(751) := X"00000000";
		ram_buffer(752) := X"00000000";
		ram_buffer(753) := X"00000000";
		ram_buffer(754) := X"00000000";
		ram_buffer(755) := X"00000000";
		ram_buffer(756) := X"00000000";
		ram_buffer(757) := X"00000000";
		ram_buffer(758) := X"00000000";
		ram_buffer(759) := X"00000000";
		ram_buffer(760) := X"00000000";
		ram_buffer(761) := X"00000000";
		ram_buffer(762) := X"00000000";
		ram_buffer(763) := X"00000000";
		ram_buffer(764) := X"00000000";
		ram_buffer(765) := X"00000000";
		ram_buffer(766) := X"00000000";
		ram_buffer(767) := X"00000000";
		ram_buffer(768) := X"00000000";
		ram_buffer(769) := X"00000000";
		ram_buffer(770) := X"00000000";
		ram_buffer(771) := X"00000000";
		ram_buffer(772) := X"00000000";
		ram_buffer(773) := X"00000000";
		ram_buffer(774) := X"00000000";
		ram_buffer(775) := X"00000000";
		ram_buffer(776) := X"00000000";
		ram_buffer(777) := X"00000000";
		ram_buffer(778) := X"00000000";
		ram_buffer(779) := X"00000000";
		ram_buffer(780) := X"00000000";
		ram_buffer(781) := X"00000000";
		ram_buffer(782) := X"00000000";
		ram_buffer(783) := X"00000000";
		ram_buffer(784) := X"00000000";
		ram_buffer(785) := X"00000000";
		ram_buffer(786) := X"00000000";
		ram_buffer(787) := X"00000000";
		ram_buffer(788) := X"00000000";
		ram_buffer(789) := X"00000000";
		ram_buffer(790) := X"00000000";
		ram_buffer(791) := X"00000000";
		ram_buffer(792) := X"00000000";
		ram_buffer(793) := X"00000000";
		ram_buffer(794) := X"00000000";
		ram_buffer(795) := X"00000000";
		ram_buffer(796) := X"00000000";
		ram_buffer(797) := X"00000000";
		ram_buffer(798) := X"00000000";
		ram_buffer(799) := X"00000000";
		ram_buffer(800) := X"00000000";
		ram_buffer(801) := X"00000000";
		ram_buffer(802) := X"00000000";
		ram_buffer(803) := X"00000000";
		ram_buffer(804) := X"00000000";
		ram_buffer(805) := X"00000000";
		ram_buffer(806) := X"00000000";
		ram_buffer(807) := X"00000000";
		ram_buffer(808) := X"00000000";
		ram_buffer(809) := X"00000000";
		ram_buffer(810) := X"00000000";
		ram_buffer(811) := X"00000000";
		ram_buffer(812) := X"00000000";
		ram_buffer(813) := X"00000000";
		ram_buffer(814) := X"00000000";
		ram_buffer(815) := X"00000000";
		ram_buffer(816) := X"00000000";
		ram_buffer(817) := X"00000000";
		ram_buffer(818) := X"00000000";
		ram_buffer(819) := X"00000000";
		ram_buffer(820) := X"00000000";
		ram_buffer(821) := X"00000000";
		ram_buffer(822) := X"00000000";
		ram_buffer(823) := X"00000000";
		ram_buffer(824) := X"00000000";
		ram_buffer(825) := X"00000000";
		ram_buffer(826) := X"00000000";
		ram_buffer(827) := X"00000000";
		ram_buffer(828) := X"00000000";
		ram_buffer(829) := X"00000000";
		ram_buffer(830) := X"00000000";
		ram_buffer(831) := X"00000000";
		ram_buffer(832) := X"00000000";
		ram_buffer(833) := X"00000000";
		ram_buffer(834) := X"00000000";
		ram_buffer(835) := X"00000000";
		ram_buffer(836) := X"00000000";
		ram_buffer(837) := X"00000000";
		ram_buffer(838) := X"00000000";
		ram_buffer(839) := X"00000000";
		ram_buffer(840) := X"00000000";
		ram_buffer(841) := X"00000000";
		ram_buffer(842) := X"00000000";
		ram_buffer(843) := X"00000000";
		ram_buffer(844) := X"00000000";
		ram_buffer(845) := X"00000000";
		ram_buffer(846) := X"00000000";
		ram_buffer(847) := X"00000000";
		ram_buffer(848) := X"00000000";
		ram_buffer(849) := X"00000000";
		ram_buffer(850) := X"00000000";
		ram_buffer(851) := X"00000000";
		ram_buffer(852) := X"00000000";
		ram_buffer(853) := X"00000000";
		ram_buffer(854) := X"00000000";
		ram_buffer(855) := X"00000000";
		ram_buffer(856) := X"00000000";
		ram_buffer(857) := X"00000000";
		ram_buffer(858) := X"00000000";
		ram_buffer(859) := X"00000000";
		ram_buffer(860) := X"00000000";
		ram_buffer(861) := X"00000000";
		ram_buffer(862) := X"00000000";
		ram_buffer(863) := X"00000000";
		ram_buffer(864) := X"00000000";
		ram_buffer(865) := X"00000000";
		ram_buffer(866) := X"00000000";
		ram_buffer(867) := X"00000000";
		ram_buffer(868) := X"00000000";
		ram_buffer(869) := X"00000000";
		ram_buffer(870) := X"00000000";
		ram_buffer(871) := X"00000000";
		ram_buffer(872) := X"00000000";
		ram_buffer(873) := X"00000000";
		ram_buffer(874) := X"00000000";
		ram_buffer(875) := X"00000000";
		ram_buffer(876) := X"00000000";
		ram_buffer(877) := X"00000000";
		ram_buffer(878) := X"00000000";
		ram_buffer(879) := X"00000000";
		ram_buffer(880) := X"00000000";
		ram_buffer(881) := X"00000000";
		ram_buffer(882) := X"00000000";
		ram_buffer(883) := X"00000000";
		ram_buffer(884) := X"00000000";
		ram_buffer(885) := X"00000000";
		ram_buffer(886) := X"00000000";
		ram_buffer(887) := X"00000000";
		ram_buffer(888) := X"00000000";
		ram_buffer(889) := X"00000000";
		ram_buffer(890) := X"00000000";
		ram_buffer(891) := X"00000000";
		ram_buffer(892) := X"00000000";
		ram_buffer(893) := X"00000000";
		ram_buffer(894) := X"00000000";
		ram_buffer(895) := X"00000000";
		ram_buffer(896) := X"00000000";
		ram_buffer(897) := X"00000000";
		ram_buffer(898) := X"00000000";
		ram_buffer(899) := X"00000000";
		ram_buffer(900) := X"00000000";
		ram_buffer(901) := X"00000000";
		ram_buffer(902) := X"00000000";
		ram_buffer(903) := X"00000000";
		ram_buffer(904) := X"00000000";
		ram_buffer(905) := X"00000000";
		ram_buffer(906) := X"00000000";
		ram_buffer(907) := X"00000000";
		ram_buffer(908) := X"00000000";
		ram_buffer(909) := X"00000000";
		ram_buffer(910) := X"00000000";
		ram_buffer(911) := X"00000000";
		ram_buffer(912) := X"00000000";
		ram_buffer(913) := X"00000000";
		ram_buffer(914) := X"00000000";
		ram_buffer(915) := X"00000000";
		ram_buffer(916) := X"00000000";
		ram_buffer(917) := X"00000000";
		ram_buffer(918) := X"00000000";
		ram_buffer(919) := X"00000000";
		ram_buffer(920) := X"00000000";
		ram_buffer(921) := X"00000000";
		ram_buffer(922) := X"00000000";
		ram_buffer(923) := X"00000000";
		ram_buffer(924) := X"00000000";
		ram_buffer(925) := X"00000000";
		ram_buffer(926) := X"00000000";
		ram_buffer(927) := X"00000000";
		ram_buffer(928) := X"00000000";
		ram_buffer(929) := X"00000000";
		ram_buffer(930) := X"00000000";
		ram_buffer(931) := X"00000000";
		ram_buffer(932) := X"00000000";
		ram_buffer(933) := X"00000000";
		ram_buffer(934) := X"00000000";
		ram_buffer(935) := X"00000000";
		ram_buffer(936) := X"00000000";
		ram_buffer(937) := X"00000000";
		ram_buffer(938) := X"00000000";
		ram_buffer(939) := X"00000000";
		ram_buffer(940) := X"00000000";
		ram_buffer(941) := X"00000000";
		ram_buffer(942) := X"00000000";
		ram_buffer(943) := X"00000000";
		ram_buffer(944) := X"00000000";
		ram_buffer(945) := X"00000000";
		ram_buffer(946) := X"00000000";
		ram_buffer(947) := X"00000000";
		ram_buffer(948) := X"00000000";
		ram_buffer(949) := X"00000000";
		ram_buffer(950) := X"00000000";
		ram_buffer(951) := X"00000000";
		ram_buffer(952) := X"00000000";
		ram_buffer(953) := X"00000000";
		ram_buffer(954) := X"00000000";
		ram_buffer(955) := X"00000000";
		ram_buffer(956) := X"00000000";
		ram_buffer(957) := X"00000000";
		ram_buffer(958) := X"00000000";
		ram_buffer(959) := X"00000000";
		ram_buffer(960) := X"00000000";
		ram_buffer(961) := X"00000000";
		ram_buffer(962) := X"00000000";
		ram_buffer(963) := X"00000000";
		ram_buffer(964) := X"00000000";
		ram_buffer(965) := X"00000000";
		ram_buffer(966) := X"00000000";
		ram_buffer(967) := X"00000000";
		ram_buffer(968) := X"00000000";
		ram_buffer(969) := X"00000000";
		ram_buffer(970) := X"00000000";
		ram_buffer(971) := X"00000000";
		ram_buffer(972) := X"00000000";
		ram_buffer(973) := X"00000000";
		ram_buffer(974) := X"00000000";
		ram_buffer(975) := X"00000000";
		ram_buffer(976) := X"00000000";
		ram_buffer(977) := X"00000000";
		ram_buffer(978) := X"00000000";
		ram_buffer(979) := X"00000000";
		ram_buffer(980) := X"00000000";
		ram_buffer(981) := X"00000000";
		ram_buffer(982) := X"00000000";
		ram_buffer(983) := X"00000000";
		ram_buffer(984) := X"00000000";
		ram_buffer(985) := X"00000000";
		ram_buffer(986) := X"00000000";
		ram_buffer(987) := X"00000000";
		ram_buffer(988) := X"00000000";
		ram_buffer(989) := X"00000000";
		ram_buffer(990) := X"00000000";
		ram_buffer(991) := X"00000000";
		ram_buffer(992) := X"00000000";
		ram_buffer(993) := X"00000000";
		ram_buffer(994) := X"00000000";
		ram_buffer(995) := X"00000000";
		ram_buffer(996) := X"00000000";
		ram_buffer(997) := X"00000000";
		ram_buffer(998) := X"00000000";
		ram_buffer(999) := X"00000000";
		ram_buffer(1000) := X"00000000";
		ram_buffer(1001) := X"00000000";
		ram_buffer(1002) := X"00000000";
		ram_buffer(1003) := X"00000000";
		ram_buffer(1004) := X"00000000";
		ram_buffer(1005) := X"00000000";
		ram_buffer(1006) := X"00000000";
		ram_buffer(1007) := X"00000000";
		ram_buffer(1008) := X"00000000";
		ram_buffer(1009) := X"00000000";
		ram_buffer(1010) := X"00000000";
		ram_buffer(1011) := X"00000000";
		ram_buffer(1012) := X"00000000";
		ram_buffer(1013) := X"00000000";
		ram_buffer(1014) := X"00000000";
		ram_buffer(1015) := X"00000000";
		ram_buffer(1016) := X"00000000";
		ram_buffer(1017) := X"00000000";
		ram_buffer(1018) := X"00000000";
		ram_buffer(1019) := X"00000000";
		ram_buffer(1020) := X"00000000";
		ram_buffer(1021) := X"00000000";
		ram_buffer(1022) := X"00000000";
		ram_buffer(1023) := X"00000000";
		ram_buffer(1024) := X"00000000";
		ram_buffer(1025) := X"00000000";
		ram_buffer(1026) := X"00000000";
		ram_buffer(1027) := X"00000000";
		ram_buffer(1028) := X"00000000";
		ram_buffer(1029) := X"00000000";
		ram_buffer(1030) := X"00000000";
		ram_buffer(1031) := X"00000000";
		ram_buffer(1032) := X"00000000";
		ram_buffer(1033) := X"00000000";
		ram_buffer(1034) := X"00000000";
		ram_buffer(1035) := X"00000000";
		ram_buffer(1036) := X"00000000";
		ram_buffer(1037) := X"00000000";
		ram_buffer(1038) := X"00000000";
		ram_buffer(1039) := X"00000000";
		ram_buffer(1040) := X"00000000";
		ram_buffer(1041) := X"00000000";
		ram_buffer(1042) := X"00000000";
		ram_buffer(1043) := X"00000000";
		ram_buffer(1044) := X"00000000";
		ram_buffer(1045) := X"00000000";
		ram_buffer(1046) := X"00000000";
		ram_buffer(1047) := X"00000000";
		ram_buffer(1048) := X"00000000";
		ram_buffer(1049) := X"00000000";
		ram_buffer(1050) := X"00000000";
		ram_buffer(1051) := X"00000000";
		ram_buffer(1052) := X"00000000";
		ram_buffer(1053) := X"00000000";
		ram_buffer(1054) := X"00000000";
		ram_buffer(1055) := X"00000000";
		ram_buffer(1056) := X"00000000";
		ram_buffer(1057) := X"00000000";
		ram_buffer(1058) := X"00000000";
		ram_buffer(1059) := X"00000000";
		ram_buffer(1060) := X"00000000";
		ram_buffer(1061) := X"00000000";
		ram_buffer(1062) := X"00000000";
		ram_buffer(1063) := X"00000000";
		ram_buffer(1064) := X"00000000";
		ram_buffer(1065) := X"00000000";
		ram_buffer(1066) := X"00000000";
		ram_buffer(1067) := X"00000000";
		ram_buffer(1068) := X"00000000";
		ram_buffer(1069) := X"00000000";
		ram_buffer(1070) := X"00000000";
		ram_buffer(1071) := X"00000000";
		ram_buffer(1072) := X"00000000";
		ram_buffer(1073) := X"00000000";
		ram_buffer(1074) := X"00000000";
		ram_buffer(1075) := X"00000000";
		ram_buffer(1076) := X"00000000";
		ram_buffer(1077) := X"00000000";
		ram_buffer(1078) := X"00000000";
		ram_buffer(1079) := X"00000000";
		ram_buffer(1080) := X"00000000";
		ram_buffer(1081) := X"00000000";
		ram_buffer(1082) := X"00000000";
		ram_buffer(1083) := X"00000000";
		ram_buffer(1084) := X"00000000";
		ram_buffer(1085) := X"00000000";
		ram_buffer(1086) := X"00000000";
		ram_buffer(1087) := X"00000000";
		ram_buffer(1088) := X"00000000";
		ram_buffer(1089) := X"00000000";
		ram_buffer(1090) := X"00000000";
		ram_buffer(1091) := X"00000000";
		ram_buffer(1092) := X"00000000";
		ram_buffer(1093) := X"00000000";
		ram_buffer(1094) := X"00000000";
		ram_buffer(1095) := X"00000000";
		ram_buffer(1096) := X"00000000";
		ram_buffer(1097) := X"00000000";
		ram_buffer(1098) := X"00000000";
		ram_buffer(1099) := X"00000000";
		ram_buffer(1100) := X"00000000";
		ram_buffer(1101) := X"00000000";
		ram_buffer(1102) := X"00000000";
		ram_buffer(1103) := X"00000000";
		ram_buffer(1104) := X"00000000";
		ram_buffer(1105) := X"00000000";
		ram_buffer(1106) := X"00000000";
		ram_buffer(1107) := X"00000000";
		ram_buffer(1108) := X"00000000";
		ram_buffer(1109) := X"00000000";
		ram_buffer(1110) := X"00000000";
		ram_buffer(1111) := X"00000000";
		ram_buffer(1112) := X"00000000";
		ram_buffer(1113) := X"00000000";
		ram_buffer(1114) := X"00000000";
		ram_buffer(1115) := X"00000000";
		ram_buffer(1116) := X"00000000";
		ram_buffer(1117) := X"00000000";
		ram_buffer(1118) := X"00000000";
		ram_buffer(1119) := X"00000000";
		ram_buffer(1120) := X"00000000";
		ram_buffer(1121) := X"00000000";
		ram_buffer(1122) := X"00000000";
		ram_buffer(1123) := X"00000000";
		ram_buffer(1124) := X"00000000";
		ram_buffer(1125) := X"00000000";
		ram_buffer(1126) := X"00000000";
		ram_buffer(1127) := X"00000000";
		ram_buffer(1128) := X"00000000";
		ram_buffer(1129) := X"00000000";
		ram_buffer(1130) := X"00000000";
		ram_buffer(1131) := X"00000000";
		ram_buffer(1132) := X"00000000";
		ram_buffer(1133) := X"00000000";
		ram_buffer(1134) := X"00000000";
		ram_buffer(1135) := X"00000000";
		ram_buffer(1136) := X"00000000";
		ram_buffer(1137) := X"00000000";
		ram_buffer(1138) := X"00000000";
		ram_buffer(1139) := X"00000000";
		ram_buffer(1140) := X"00000000";
		ram_buffer(1141) := X"00000000";
		ram_buffer(1142) := X"00000000";
		ram_buffer(1143) := X"00000000";
		ram_buffer(1144) := X"00000000";
		ram_buffer(1145) := X"00000000";
		ram_buffer(1146) := X"00000000";
		ram_buffer(1147) := X"00000000";
		ram_buffer(1148) := X"00000000";
		ram_buffer(1149) := X"00000000";
		ram_buffer(1150) := X"00000000";
		ram_buffer(1151) := X"00000000";
		ram_buffer(1152) := X"00000000";
		ram_buffer(1153) := X"00000000";
		ram_buffer(1154) := X"00000000";
		ram_buffer(1155) := X"00000000";
		ram_buffer(1156) := X"00000000";
		ram_buffer(1157) := X"00000000";
		ram_buffer(1158) := X"00000000";
		ram_buffer(1159) := X"00000000";
		ram_buffer(1160) := X"00000000";
		ram_buffer(1161) := X"00000000";
		ram_buffer(1162) := X"00000000";
		ram_buffer(1163) := X"00000000";
		ram_buffer(1164) := X"00000000";
		ram_buffer(1165) := X"00000000";
		ram_buffer(1166) := X"00000000";
		ram_buffer(1167) := X"00000000";
		ram_buffer(1168) := X"00000000";
		ram_buffer(1169) := X"00000000";
		ram_buffer(1170) := X"00000000";
		ram_buffer(1171) := X"00000000";
		ram_buffer(1172) := X"00000000";
		ram_buffer(1173) := X"00000000";
		ram_buffer(1174) := X"00000000";
		ram_buffer(1175) := X"00000000";
		ram_buffer(1176) := X"00000000";
		ram_buffer(1177) := X"00000000";
		ram_buffer(1178) := X"00000000";
		ram_buffer(1179) := X"00000000";
		ram_buffer(1180) := X"00000000";
		ram_buffer(1181) := X"00000000";
		ram_buffer(1182) := X"00000000";
		ram_buffer(1183) := X"00000000";
		ram_buffer(1184) := X"00000000";
		ram_buffer(1185) := X"00000000";
		ram_buffer(1186) := X"00000000";
		ram_buffer(1187) := X"00000000";
		ram_buffer(1188) := X"00000000";
		ram_buffer(1189) := X"00000000";
		ram_buffer(1190) := X"00000000";
		ram_buffer(1191) := X"00000000";
		ram_buffer(1192) := X"00000000";
		ram_buffer(1193) := X"00000000";
		ram_buffer(1194) := X"00000000";
		ram_buffer(1195) := X"00000000";
		ram_buffer(1196) := X"00000000";
		ram_buffer(1197) := X"00000000";
		ram_buffer(1198) := X"00000000";
		ram_buffer(1199) := X"00000000";
		ram_buffer(1200) := X"00000000";
		ram_buffer(1201) := X"00000000";
		ram_buffer(1202) := X"00000000";
		ram_buffer(1203) := X"00000000";
		ram_buffer(1204) := X"00000000";
		ram_buffer(1205) := X"00000000";
		ram_buffer(1206) := X"00000000";
		ram_buffer(1207) := X"00000000";
		ram_buffer(1208) := X"00000000";
		ram_buffer(1209) := X"00000000";
		ram_buffer(1210) := X"00000000";
		ram_buffer(1211) := X"00000000";
		ram_buffer(1212) := X"00000000";
		ram_buffer(1213) := X"00000000";
		ram_buffer(1214) := X"00000000";
		ram_buffer(1215) := X"00000000";
		ram_buffer(1216) := X"00000000";
		ram_buffer(1217) := X"00000000";
		ram_buffer(1218) := X"00000000";
		ram_buffer(1219) := X"00000000";
		ram_buffer(1220) := X"00000000";
		ram_buffer(1221) := X"00000000";
		ram_buffer(1222) := X"00000000";
		ram_buffer(1223) := X"00000000";
		ram_buffer(1224) := X"00000000";
		ram_buffer(1225) := X"00000000";
		ram_buffer(1226) := X"00000000";
		ram_buffer(1227) := X"00000000";
		ram_buffer(1228) := X"00000000";
		ram_buffer(1229) := X"00000000";
		ram_buffer(1230) := X"00000000";
		ram_buffer(1231) := X"00000000";
		ram_buffer(1232) := X"00000000";
		ram_buffer(1233) := X"00000000";
		ram_buffer(1234) := X"00000000";
		ram_buffer(1235) := X"00000000";
		ram_buffer(1236) := X"00000000";
		ram_buffer(1237) := X"00000000";
		ram_buffer(1238) := X"00000000";
		ram_buffer(1239) := X"00000000";
		ram_buffer(1240) := X"00000000";
		ram_buffer(1241) := X"00000000";
		ram_buffer(1242) := X"00000000";
		ram_buffer(1243) := X"00000000";
		ram_buffer(1244) := X"00000000";
		ram_buffer(1245) := X"00000000";
		ram_buffer(1246) := X"00000000";
		ram_buffer(1247) := X"00000000";
		ram_buffer(1248) := X"00000000";
		ram_buffer(1249) := X"00000000";
		ram_buffer(1250) := X"00000000";
		ram_buffer(1251) := X"00000000";
		ram_buffer(1252) := X"00000000";
		ram_buffer(1253) := X"00000000";
		ram_buffer(1254) := X"00000000";
		ram_buffer(1255) := X"00000000";
		ram_buffer(1256) := X"00000000";
		ram_buffer(1257) := X"00000000";
		ram_buffer(1258) := X"00000000";
		ram_buffer(1259) := X"00000000";
		ram_buffer(1260) := X"00000000";
		ram_buffer(1261) := X"00000000";
		ram_buffer(1262) := X"00000000";
		ram_buffer(1263) := X"00000000";
		ram_buffer(1264) := X"00000000";
		ram_buffer(1265) := X"00000000";
		ram_buffer(1266) := X"00000000";
		ram_buffer(1267) := X"00000000";
		ram_buffer(1268) := X"00000000";
		ram_buffer(1269) := X"00000000";
		ram_buffer(1270) := X"00000000";
		ram_buffer(1271) := X"00000000";
		ram_buffer(1272) := X"00000000";
		ram_buffer(1273) := X"00000000";
		ram_buffer(1274) := X"00000000";
		ram_buffer(1275) := X"00000000";
		ram_buffer(1276) := X"00000000";
		ram_buffer(1277) := X"00000000";
		ram_buffer(1278) := X"00000000";
		ram_buffer(1279) := X"00000000";
		ram_buffer(1280) := X"00000000";
		ram_buffer(1281) := X"00000000";
		ram_buffer(1282) := X"00000000";
		ram_buffer(1283) := X"00000000";
		ram_buffer(1284) := X"00000000";
		ram_buffer(1285) := X"00000000";
		ram_buffer(1286) := X"00000000";
		ram_buffer(1287) := X"00000000";
		ram_buffer(1288) := X"00000000";
		ram_buffer(1289) := X"00000000";
		ram_buffer(1290) := X"00000000";
		ram_buffer(1291) := X"00000000";
		ram_buffer(1292) := X"00000000";
		ram_buffer(1293) := X"00000000";
		ram_buffer(1294) := X"00000000";
		ram_buffer(1295) := X"00000000";
		ram_buffer(1296) := X"00000000";
		ram_buffer(1297) := X"00000000";
		ram_buffer(1298) := X"00000000";
		ram_buffer(1299) := X"00000000";
		ram_buffer(1300) := X"00000000";
		ram_buffer(1301) := X"00000000";
		ram_buffer(1302) := X"00000000";
		ram_buffer(1303) := X"00000000";
		ram_buffer(1304) := X"00000000";
		ram_buffer(1305) := X"00000000";
		ram_buffer(1306) := X"00000000";
		ram_buffer(1307) := X"00000000";
		ram_buffer(1308) := X"00000000";
		ram_buffer(1309) := X"00000000";
		ram_buffer(1310) := X"00000000";
		ram_buffer(1311) := X"00000000";
		ram_buffer(1312) := X"00000000";
		ram_buffer(1313) := X"00000000";
		ram_buffer(1314) := X"00000000";
		ram_buffer(1315) := X"00000000";
		ram_buffer(1316) := X"00000000";
		ram_buffer(1317) := X"00000000";
		ram_buffer(1318) := X"00000000";
		ram_buffer(1319) := X"00000000";
		ram_buffer(1320) := X"00000000";
		ram_buffer(1321) := X"00000000";
		ram_buffer(1322) := X"00000000";
		ram_buffer(1323) := X"00000000";
		ram_buffer(1324) := X"00000000";
		ram_buffer(1325) := X"00000000";
		ram_buffer(1326) := X"00000000";
		ram_buffer(1327) := X"00000000";
		ram_buffer(1328) := X"00000000";
		ram_buffer(1329) := X"00000000";
		ram_buffer(1330) := X"00000000";
		ram_buffer(1331) := X"00000000";
		ram_buffer(1332) := X"00000000";
		ram_buffer(1333) := X"00000000";
		ram_buffer(1334) := X"00000000";
		ram_buffer(1335) := X"00000000";
		ram_buffer(1336) := X"00000000";
		ram_buffer(1337) := X"00000000";
		ram_buffer(1338) := X"00000000";
		ram_buffer(1339) := X"00000000";
		ram_buffer(1340) := X"00000000";
		ram_buffer(1341) := X"00000000";
		ram_buffer(1342) := X"00000000";
		ram_buffer(1343) := X"00000000";
		ram_buffer(1344) := X"00000000";
		ram_buffer(1345) := X"00000000";
		ram_buffer(1346) := X"00000000";
		ram_buffer(1347) := X"00000000";
		ram_buffer(1348) := X"00000000";
		ram_buffer(1349) := X"00000000";
		ram_buffer(1350) := X"00000000";
		ram_buffer(1351) := X"00000000";
		ram_buffer(1352) := X"00000000";
		ram_buffer(1353) := X"00000000";
		ram_buffer(1354) := X"00000000";
		ram_buffer(1355) := X"00000000";
		ram_buffer(1356) := X"00000000";
		ram_buffer(1357) := X"00000000";
		ram_buffer(1358) := X"00000000";
		ram_buffer(1359) := X"00000000";
		ram_buffer(1360) := X"00000000";
		ram_buffer(1361) := X"00000000";
		ram_buffer(1362) := X"00000000";
		ram_buffer(1363) := X"00000000";
		ram_buffer(1364) := X"00000000";
		ram_buffer(1365) := X"00000000";
		ram_buffer(1366) := X"00000000";
		ram_buffer(1367) := X"00000000";
		ram_buffer(1368) := X"00000000";
		ram_buffer(1369) := X"00000000";
		ram_buffer(1370) := X"00000000";
		ram_buffer(1371) := X"00000000";
		ram_buffer(1372) := X"00000000";
		ram_buffer(1373) := X"00000000";
		ram_buffer(1374) := X"00000000";
		ram_buffer(1375) := X"00000000";
		ram_buffer(1376) := X"00000000";
		ram_buffer(1377) := X"00000000";
		ram_buffer(1378) := X"00000000";
		ram_buffer(1379) := X"00000000";
		ram_buffer(1380) := X"00000000";
		ram_buffer(1381) := X"00000000";
		ram_buffer(1382) := X"00000000";
		ram_buffer(1383) := X"00000000";
		ram_buffer(1384) := X"00000000";
		ram_buffer(1385) := X"00000000";
		ram_buffer(1386) := X"00000000";
		ram_buffer(1387) := X"00000000";
		ram_buffer(1388) := X"00000000";
		ram_buffer(1389) := X"00000000";
		ram_buffer(1390) := X"00000000";
		ram_buffer(1391) := X"00000000";
		ram_buffer(1392) := X"00000000";
		ram_buffer(1393) := X"00000000";
		ram_buffer(1394) := X"00000000";
		ram_buffer(1395) := X"00000000";
		ram_buffer(1396) := X"00000000";
		ram_buffer(1397) := X"00000000";
		ram_buffer(1398) := X"00000000";
		ram_buffer(1399) := X"00000000";
		ram_buffer(1400) := X"00000000";
		ram_buffer(1401) := X"00000000";
		ram_buffer(1402) := X"00000000";
		ram_buffer(1403) := X"00000000";
		ram_buffer(1404) := X"00000000";
		ram_buffer(1405) := X"00000000";
		ram_buffer(1406) := X"00000000";
		ram_buffer(1407) := X"00000000";
		ram_buffer(1408) := X"00000000";
		ram_buffer(1409) := X"00000000";
		ram_buffer(1410) := X"00000000";
		ram_buffer(1411) := X"00000000";
		ram_buffer(1412) := X"00000000";
		ram_buffer(1413) := X"00000000";
		ram_buffer(1414) := X"00000000";
		ram_buffer(1415) := X"00000000";
		ram_buffer(1416) := X"00000000";
		ram_buffer(1417) := X"00000000";
		ram_buffer(1418) := X"00000000";
		ram_buffer(1419) := X"00000000";
		ram_buffer(1420) := X"00000000";
		ram_buffer(1421) := X"00000000";
		ram_buffer(1422) := X"00000000";
		ram_buffer(1423) := X"00000000";
		ram_buffer(1424) := X"00000000";
		ram_buffer(1425) := X"00000000";
		ram_buffer(1426) := X"00000000";
		ram_buffer(1427) := X"00000000";
		ram_buffer(1428) := X"00000000";
		ram_buffer(1429) := X"00000000";
		ram_buffer(1430) := X"00000000";
		ram_buffer(1431) := X"00000000";
		ram_buffer(1432) := X"00000000";
		ram_buffer(1433) := X"00000000";
		ram_buffer(1434) := X"00000000";
		ram_buffer(1435) := X"00000000";
		ram_buffer(1436) := X"00000000";
		ram_buffer(1437) := X"00000000";
		ram_buffer(1438) := X"00000000";
		ram_buffer(1439) := X"00000000";
		ram_buffer(1440) := X"00000000";
		ram_buffer(1441) := X"00000000";
		ram_buffer(1442) := X"00000000";
		ram_buffer(1443) := X"00000000";
		ram_buffer(1444) := X"00000000";
		ram_buffer(1445) := X"00000000";
		ram_buffer(1446) := X"00000000";
		ram_buffer(1447) := X"00000000";
		ram_buffer(1448) := X"00000000";
		ram_buffer(1449) := X"00000000";
		ram_buffer(1450) := X"00000000";
		ram_buffer(1451) := X"00000000";
		ram_buffer(1452) := X"00000000";
		ram_buffer(1453) := X"00000000";
		ram_buffer(1454) := X"00000000";
		ram_buffer(1455) := X"00000000";
		ram_buffer(1456) := X"00000000";
		ram_buffer(1457) := X"00000000";
		ram_buffer(1458) := X"00000000";
		ram_buffer(1459) := X"00000000";
		ram_buffer(1460) := X"00000000";
		ram_buffer(1461) := X"00000000";
		ram_buffer(1462) := X"00000000";
		ram_buffer(1463) := X"00000000";
		ram_buffer(1464) := X"00000000";
		ram_buffer(1465) := X"00000000";
		ram_buffer(1466) := X"00000000";
		ram_buffer(1467) := X"00000000";
		ram_buffer(1468) := X"00000000";
		ram_buffer(1469) := X"00000000";
		ram_buffer(1470) := X"00000000";
		ram_buffer(1471) := X"00000000";
		ram_buffer(1472) := X"00000000";
		ram_buffer(1473) := X"00000000";
		ram_buffer(1474) := X"00000000";
		ram_buffer(1475) := X"00000000";
		ram_buffer(1476) := X"00000000";
		ram_buffer(1477) := X"00000000";
		ram_buffer(1478) := X"00000000";
		ram_buffer(1479) := X"00000000";
		ram_buffer(1480) := X"00000000";
		ram_buffer(1481) := X"00000000";
		ram_buffer(1482) := X"00000000";
		ram_buffer(1483) := X"00000000";
		ram_buffer(1484) := X"00000000";
		ram_buffer(1485) := X"00000000";
		ram_buffer(1486) := X"00000000";
		ram_buffer(1487) := X"00000000";
		ram_buffer(1488) := X"00000000";
		ram_buffer(1489) := X"00000000";
		ram_buffer(1490) := X"00000000";
		ram_buffer(1491) := X"00000000";
		ram_buffer(1492) := X"00000000";
		ram_buffer(1493) := X"00000000";
		ram_buffer(1494) := X"00000000";
		ram_buffer(1495) := X"00000000";
		ram_buffer(1496) := X"00000000";
		ram_buffer(1497) := X"00000000";
		ram_buffer(1498) := X"00000000";
		ram_buffer(1499) := X"00000000";
		ram_buffer(1500) := X"00000000";
		ram_buffer(1501) := X"00000000";
		ram_buffer(1502) := X"00000000";
		ram_buffer(1503) := X"00000000";
		ram_buffer(1504) := X"00000000";
		ram_buffer(1505) := X"00000000";
		ram_buffer(1506) := X"00000000";
		ram_buffer(1507) := X"00000000";
		ram_buffer(1508) := X"00000000";
		ram_buffer(1509) := X"00000000";
		ram_buffer(1510) := X"00000000";
		ram_buffer(1511) := X"00000000";
		ram_buffer(1512) := X"00000000";
		ram_buffer(1513) := X"00000000";
		ram_buffer(1514) := X"00000000";
		ram_buffer(1515) := X"00000000";
		ram_buffer(1516) := X"00000000";
		ram_buffer(1517) := X"00000000";
		ram_buffer(1518) := X"00000000";
		ram_buffer(1519) := X"00000000";
		ram_buffer(1520) := X"00000000";
		ram_buffer(1521) := X"00000000";
		ram_buffer(1522) := X"00000000";
		ram_buffer(1523) := X"00000000";
		ram_buffer(1524) := X"00000000";
		ram_buffer(1525) := X"00000000";
		ram_buffer(1526) := X"00000000";
		ram_buffer(1527) := X"00000000";
		ram_buffer(1528) := X"00000000";
		ram_buffer(1529) := X"00000000";
		ram_buffer(1530) := X"00000000";
		ram_buffer(1531) := X"00000000";
		ram_buffer(1532) := X"00000000";
		ram_buffer(1533) := X"00000000";
		ram_buffer(1534) := X"00000000";
		ram_buffer(1535) := X"00000000";
		ram_buffer(1536) := X"00000000";
		ram_buffer(1537) := X"00000000";
		ram_buffer(1538) := X"00000000";
		ram_buffer(1539) := X"00000000";
		ram_buffer(1540) := X"00000000";
		ram_buffer(1541) := X"00000000";
		ram_buffer(1542) := X"00000000";
		ram_buffer(1543) := X"00000000";
		ram_buffer(1544) := X"00000000";
		ram_buffer(1545) := X"00000000";
		ram_buffer(1546) := X"00000000";
		ram_buffer(1547) := X"00000000";
		ram_buffer(1548) := X"00000000";
		ram_buffer(1549) := X"00000000";
		ram_buffer(1550) := X"00000000";
		ram_buffer(1551) := X"00000000";
		ram_buffer(1552) := X"00000000";
		ram_buffer(1553) := X"00000000";
		ram_buffer(1554) := X"00000000";
		ram_buffer(1555) := X"00000000";
		ram_buffer(1556) := X"00000000";
		ram_buffer(1557) := X"00000000";
		ram_buffer(1558) := X"00000000";
		ram_buffer(1559) := X"00000000";
		ram_buffer(1560) := X"00000000";
		ram_buffer(1561) := X"00000000";
		ram_buffer(1562) := X"00000000";
		ram_buffer(1563) := X"00000000";
		ram_buffer(1564) := X"00000000";
		ram_buffer(1565) := X"00000000";
		ram_buffer(1566) := X"00000000";
		ram_buffer(1567) := X"00000000";
		ram_buffer(1568) := X"00000000";
		ram_buffer(1569) := X"00000000";
		ram_buffer(1570) := X"00000000";
		ram_buffer(1571) := X"00000000";
		ram_buffer(1572) := X"00000000";
		ram_buffer(1573) := X"00000000";
		ram_buffer(1574) := X"00000000";
		ram_buffer(1575) := X"00000000";
		ram_buffer(1576) := X"00000000";
		ram_buffer(1577) := X"00000000";
		ram_buffer(1578) := X"00000000";
		ram_buffer(1579) := X"00000000";
		ram_buffer(1580) := X"00000000";
		ram_buffer(1581) := X"00000000";
		ram_buffer(1582) := X"00000000";
		ram_buffer(1583) := X"00000000";
		ram_buffer(1584) := X"00000000";
		ram_buffer(1585) := X"00000000";
		ram_buffer(1586) := X"00000000";
		ram_buffer(1587) := X"00000000";
		ram_buffer(1588) := X"00000000";
		ram_buffer(1589) := X"00000000";
		ram_buffer(1590) := X"00000000";
		ram_buffer(1591) := X"00000000";
		ram_buffer(1592) := X"00000000";
		ram_buffer(1593) := X"00000000";
		ram_buffer(1594) := X"00000000";
		ram_buffer(1595) := X"00000000";
		ram_buffer(1596) := X"00000000";
		ram_buffer(1597) := X"00000000";
		ram_buffer(1598) := X"00000000";
		ram_buffer(1599) := X"00000000";
		ram_buffer(1600) := X"00000000";
		ram_buffer(1601) := X"00000000";
		ram_buffer(1602) := X"00000000";
		ram_buffer(1603) := X"00000000";
		ram_buffer(1604) := X"00000000";
		ram_buffer(1605) := X"00000000";
		ram_buffer(1606) := X"00000000";
		ram_buffer(1607) := X"00000000";
		ram_buffer(1608) := X"00000000";
		ram_buffer(1609) := X"00000000";
		ram_buffer(1610) := X"00000000";
		ram_buffer(1611) := X"00000000";
		ram_buffer(1612) := X"00000000";
		ram_buffer(1613) := X"00000000";
		ram_buffer(1614) := X"00000000";
		ram_buffer(1615) := X"00000000";
		ram_buffer(1616) := X"00000000";
		ram_buffer(1617) := X"00000000";
		ram_buffer(1618) := X"00000000";
		ram_buffer(1619) := X"00000000";
		ram_buffer(1620) := X"00000000";
		ram_buffer(1621) := X"00000000";
		ram_buffer(1622) := X"00000000";
		ram_buffer(1623) := X"00000000";
		ram_buffer(1624) := X"00000000";
		ram_buffer(1625) := X"00000000";
		ram_buffer(1626) := X"00000000";
		ram_buffer(1627) := X"00000000";
		ram_buffer(1628) := X"00000000";
		ram_buffer(1629) := X"00000000";
		ram_buffer(1630) := X"00000000";
		ram_buffer(1631) := X"00000000";
		ram_buffer(1632) := X"00000000";
		ram_buffer(1633) := X"00000000";
		ram_buffer(1634) := X"00000000";
		ram_buffer(1635) := X"00000000";
		ram_buffer(1636) := X"00000000";
		ram_buffer(1637) := X"00000000";
		ram_buffer(1638) := X"00000000";
		ram_buffer(1639) := X"00000000";
		ram_buffer(1640) := X"00000000";
		ram_buffer(1641) := X"00000000";
		ram_buffer(1642) := X"00000000";
		ram_buffer(1643) := X"00000000";
		ram_buffer(1644) := X"00000000";
		ram_buffer(1645) := X"00000000";
		ram_buffer(1646) := X"00000000";
		ram_buffer(1647) := X"00000000";
		ram_buffer(1648) := X"00000000";
		ram_buffer(1649) := X"00000000";
		ram_buffer(1650) := X"00000000";
		ram_buffer(1651) := X"00000000";
		ram_buffer(1652) := X"00000000";
		ram_buffer(1653) := X"00000000";
		ram_buffer(1654) := X"00000000";
		ram_buffer(1655) := X"00000000";
		ram_buffer(1656) := X"00000000";
		ram_buffer(1657) := X"00000000";
		ram_buffer(1658) := X"00000000";
		ram_buffer(1659) := X"00000000";
		ram_buffer(1660) := X"00000000";
		ram_buffer(1661) := X"00000000";
		ram_buffer(1662) := X"00000000";
		ram_buffer(1663) := X"00000000";
		ram_buffer(1664) := X"00000000";
		ram_buffer(1665) := X"00000000";
		ram_buffer(1666) := X"00000000";
		ram_buffer(1667) := X"00000000";
		ram_buffer(1668) := X"00000000";
		ram_buffer(1669) := X"00000000";
		ram_buffer(1670) := X"00000000";
		ram_buffer(1671) := X"00000000";
		ram_buffer(1672) := X"00000000";
		ram_buffer(1673) := X"00000000";
		ram_buffer(1674) := X"00000000";
		ram_buffer(1675) := X"00000000";
		ram_buffer(1676) := X"00000000";
		ram_buffer(1677) := X"00000000";
		ram_buffer(1678) := X"00000000";
		ram_buffer(1679) := X"00000000";
		ram_buffer(1680) := X"00000000";
		ram_buffer(1681) := X"00000000";
		ram_buffer(1682) := X"00000000";
		ram_buffer(1683) := X"00000000";
		ram_buffer(1684) := X"00000000";
		ram_buffer(1685) := X"00000000";
		ram_buffer(1686) := X"00000000";
		ram_buffer(1687) := X"00000000";
		ram_buffer(1688) := X"00000000";
		ram_buffer(1689) := X"00000000";
		ram_buffer(1690) := X"00000000";
		ram_buffer(1691) := X"00000000";
		ram_buffer(1692) := X"00000000";
		ram_buffer(1693) := X"00000000";
		ram_buffer(1694) := X"00000000";
		ram_buffer(1695) := X"00000000";
		ram_buffer(1696) := X"00000000";
		ram_buffer(1697) := X"00000000";
		ram_buffer(1698) := X"00000000";
		ram_buffer(1699) := X"00000000";
		ram_buffer(1700) := X"00000000";
		ram_buffer(1701) := X"00000000";
		ram_buffer(1702) := X"00000000";
		ram_buffer(1703) := X"00000000";
		ram_buffer(1704) := X"00000000";
		ram_buffer(1705) := X"00000000";
		ram_buffer(1706) := X"00000000";
		ram_buffer(1707) := X"00000000";
		ram_buffer(1708) := X"00000000";
		ram_buffer(1709) := X"00000000";
		ram_buffer(1710) := X"00000000";
		ram_buffer(1711) := X"00000000";
		ram_buffer(1712) := X"00000000";
		ram_buffer(1713) := X"00000000";
		ram_buffer(1714) := X"00000000";
		ram_buffer(1715) := X"00000000";
		ram_buffer(1716) := X"00000000";
		ram_buffer(1717) := X"00000000";
		ram_buffer(1718) := X"00000000";
		ram_buffer(1719) := X"00000000";
		ram_buffer(1720) := X"00000000";
		ram_buffer(1721) := X"00000000";
		ram_buffer(1722) := X"00000000";
		ram_buffer(1723) := X"00000000";
		ram_buffer(1724) := X"00000000";
		ram_buffer(1725) := X"00000000";
		ram_buffer(1726) := X"00000000";
		ram_buffer(1727) := X"00000000";
		ram_buffer(1728) := X"00000000";
		ram_buffer(1729) := X"00000000";
		ram_buffer(1730) := X"00000000";
		ram_buffer(1731) := X"00000000";
		ram_buffer(1732) := X"00000000";
		ram_buffer(1733) := X"00000000";
		ram_buffer(1734) := X"00000000";
		ram_buffer(1735) := X"00000000";
		ram_buffer(1736) := X"00000000";
		ram_buffer(1737) := X"00000000";
		ram_buffer(1738) := X"00000000";
		ram_buffer(1739) := X"00000000";
		ram_buffer(1740) := X"00000000";
		ram_buffer(1741) := X"00000000";
		ram_buffer(1742) := X"00000000";
		ram_buffer(1743) := X"00000000";
		ram_buffer(1744) := X"00000000";
		ram_buffer(1745) := X"00000000";
		ram_buffer(1746) := X"00000000";
		ram_buffer(1747) := X"00000000";
		ram_buffer(1748) := X"00000000";
		ram_buffer(1749) := X"00000000";
		ram_buffer(1750) := X"00000000";
		ram_buffer(1751) := X"00000000";
		ram_buffer(1752) := X"00000000";
		ram_buffer(1753) := X"00000000";
		ram_buffer(1754) := X"00000000";
		ram_buffer(1755) := X"00000000";
		ram_buffer(1756) := X"00000000";
		ram_buffer(1757) := X"00000000";
		ram_buffer(1758) := X"00000000";
		ram_buffer(1759) := X"00000000";
		ram_buffer(1760) := X"00000000";
		ram_buffer(1761) := X"00000000";
		ram_buffer(1762) := X"00000000";
		ram_buffer(1763) := X"00000000";
		ram_buffer(1764) := X"00000000";
		ram_buffer(1765) := X"00000000";
		ram_buffer(1766) := X"00000000";
		ram_buffer(1767) := X"00000000";
		ram_buffer(1768) := X"00000000";
		ram_buffer(1769) := X"00000000";
		ram_buffer(1770) := X"00000000";
		ram_buffer(1771) := X"00000000";
		ram_buffer(1772) := X"00000000";
		ram_buffer(1773) := X"00000000";
		ram_buffer(1774) := X"00000000";
		ram_buffer(1775) := X"00000000";
		ram_buffer(1776) := X"00000000";
		ram_buffer(1777) := X"00000000";
		ram_buffer(1778) := X"00000000";
		ram_buffer(1779) := X"00000000";
		ram_buffer(1780) := X"00000000";
		ram_buffer(1781) := X"00000000";
		ram_buffer(1782) := X"00000000";
		ram_buffer(1783) := X"00000000";
		ram_buffer(1784) := X"00000000";
		ram_buffer(1785) := X"00000000";
		ram_buffer(1786) := X"00000000";
		ram_buffer(1787) := X"00000000";
		ram_buffer(1788) := X"00000000";
		ram_buffer(1789) := X"00000000";
		ram_buffer(1790) := X"00000000";
		ram_buffer(1791) := X"00000000";
		ram_buffer(1792) := X"00000000";
		ram_buffer(1793) := X"00000000";
		ram_buffer(1794) := X"00000000";
		ram_buffer(1795) := X"00000000";
		ram_buffer(1796) := X"00000000";
		ram_buffer(1797) := X"00000000";
		ram_buffer(1798) := X"00000000";
		ram_buffer(1799) := X"00000000";
		ram_buffer(1800) := X"00000000";
		ram_buffer(1801) := X"00000000";
		ram_buffer(1802) := X"00000000";
		ram_buffer(1803) := X"00000000";
		ram_buffer(1804) := X"00000000";
		ram_buffer(1805) := X"00000000";
		ram_buffer(1806) := X"00000000";
		ram_buffer(1807) := X"00000000";
		ram_buffer(1808) := X"00000000";
		ram_buffer(1809) := X"00000000";
		ram_buffer(1810) := X"00000000";
		ram_buffer(1811) := X"00000000";
		ram_buffer(1812) := X"00000000";
		ram_buffer(1813) := X"00000000";
		ram_buffer(1814) := X"00000000";
		ram_buffer(1815) := X"00000000";
		ram_buffer(1816) := X"00000000";
		ram_buffer(1817) := X"00000000";
		ram_buffer(1818) := X"00000000";
		ram_buffer(1819) := X"00000000";
		ram_buffer(1820) := X"00000000";
		ram_buffer(1821) := X"00000000";
		ram_buffer(1822) := X"00000000";
		ram_buffer(1823) := X"00000000";
		ram_buffer(1824) := X"00000000";
		ram_buffer(1825) := X"00000000";
		ram_buffer(1826) := X"00000000";
		ram_buffer(1827) := X"00000000";
		ram_buffer(1828) := X"00000000";
		ram_buffer(1829) := X"00000000";
		ram_buffer(1830) := X"00000000";
		ram_buffer(1831) := X"00000000";
		ram_buffer(1832) := X"00000000";
		ram_buffer(1833) := X"00000000";
		ram_buffer(1834) := X"00000000";
		ram_buffer(1835) := X"00000000";
		ram_buffer(1836) := X"00000000";
		ram_buffer(1837) := X"00000000";
		ram_buffer(1838) := X"00000000";
		ram_buffer(1839) := X"00000000";
		ram_buffer(1840) := X"00000000";
		ram_buffer(1841) := X"00000000";
		ram_buffer(1842) := X"00000000";
		ram_buffer(1843) := X"00000000";
		ram_buffer(1844) := X"00000000";
		ram_buffer(1845) := X"00000000";
		ram_buffer(1846) := X"00000000";
		ram_buffer(1847) := X"00000000";
		ram_buffer(1848) := X"00000000";
		ram_buffer(1849) := X"00000000";
		ram_buffer(1850) := X"00000000";
		ram_buffer(1851) := X"00000000";
		ram_buffer(1852) := X"00000000";
		ram_buffer(1853) := X"00000000";
		ram_buffer(1854) := X"00000000";
		ram_buffer(1855) := X"00000000";
		ram_buffer(1856) := X"00000000";
		ram_buffer(1857) := X"00000000";
		ram_buffer(1858) := X"00000000";
		ram_buffer(1859) := X"00000000";
		ram_buffer(1860) := X"00000000";
		ram_buffer(1861) := X"00000000";
		ram_buffer(1862) := X"00000000";
		ram_buffer(1863) := X"00000000";
		ram_buffer(1864) := X"00000000";
		ram_buffer(1865) := X"00000000";
		ram_buffer(1866) := X"00000000";
		ram_buffer(1867) := X"00000000";
		ram_buffer(1868) := X"00000000";
		ram_buffer(1869) := X"00000000";
		ram_buffer(1870) := X"00000000";
		ram_buffer(1871) := X"00000000";
		ram_buffer(1872) := X"00000000";
		ram_buffer(1873) := X"00000000";
		ram_buffer(1874) := X"00000000";
		ram_buffer(1875) := X"00000000";
		ram_buffer(1876) := X"00000000";
		ram_buffer(1877) := X"00000000";
		ram_buffer(1878) := X"00000000";
		ram_buffer(1879) := X"00000000";
		ram_buffer(1880) := X"00000000";
		ram_buffer(1881) := X"00000000";
		ram_buffer(1882) := X"00000000";
		ram_buffer(1883) := X"00000000";
		ram_buffer(1884) := X"00000000";
		ram_buffer(1885) := X"00000000";
		ram_buffer(1886) := X"00000000";
		ram_buffer(1887) := X"00000000";
		ram_buffer(1888) := X"00000000";
		ram_buffer(1889) := X"00000000";
		ram_buffer(1890) := X"00000000";
		ram_buffer(1891) := X"00000000";
		ram_buffer(1892) := X"00000000";
		ram_buffer(1893) := X"00000000";
		ram_buffer(1894) := X"00000000";
		ram_buffer(1895) := X"00000000";
		ram_buffer(1896) := X"00000000";
		ram_buffer(1897) := X"00000000";
		ram_buffer(1898) := X"00000000";
		ram_buffer(1899) := X"00000000";
		ram_buffer(1900) := X"00000000";
		ram_buffer(1901) := X"00000000";
		ram_buffer(1902) := X"00000000";
		ram_buffer(1903) := X"00000000";
		ram_buffer(1904) := X"00000000";
		ram_buffer(1905) := X"00000000";
		ram_buffer(1906) := X"00000000";
		ram_buffer(1907) := X"00000000";
		ram_buffer(1908) := X"00000000";
		ram_buffer(1909) := X"00000000";
		ram_buffer(1910) := X"00000000";
		ram_buffer(1911) := X"00000000";
		ram_buffer(1912) := X"00000000";
		ram_buffer(1913) := X"00000000";
		ram_buffer(1914) := X"00000000";
		ram_buffer(1915) := X"00000000";
		ram_buffer(1916) := X"00000000";
		ram_buffer(1917) := X"00000000";
		ram_buffer(1918) := X"00000000";
		ram_buffer(1919) := X"00000000";
		ram_buffer(1920) := X"00000000";
		ram_buffer(1921) := X"00000000";
		ram_buffer(1922) := X"00000000";
		ram_buffer(1923) := X"00000000";
		ram_buffer(1924) := X"00000000";
		ram_buffer(1925) := X"00000000";
		ram_buffer(1926) := X"00000000";
		ram_buffer(1927) := X"00000000";
		ram_buffer(1928) := X"00000000";
		ram_buffer(1929) := X"00000000";
		ram_buffer(1930) := X"00000000";
		ram_buffer(1931) := X"00000000";
		ram_buffer(1932) := X"00000000";
		ram_buffer(1933) := X"00000000";
		ram_buffer(1934) := X"00000000";
		ram_buffer(1935) := X"00000000";
		ram_buffer(1936) := X"00000000";
		ram_buffer(1937) := X"00000000";
		ram_buffer(1938) := X"00000000";
		ram_buffer(1939) := X"00000000";
		ram_buffer(1940) := X"00000000";
		ram_buffer(1941) := X"00000000";
		ram_buffer(1942) := X"00000000";
		ram_buffer(1943) := X"00000000";
		ram_buffer(1944) := X"00000000";
		ram_buffer(1945) := X"00000000";
		ram_buffer(1946) := X"00000000";
		ram_buffer(1947) := X"00000000";
		ram_buffer(1948) := X"00000000";
		ram_buffer(1949) := X"00000000";
		ram_buffer(1950) := X"00000000";
		ram_buffer(1951) := X"00000000";
		ram_buffer(1952) := X"00000000";
		ram_buffer(1953) := X"00000000";
		ram_buffer(1954) := X"00000000";
		ram_buffer(1955) := X"00000000";
		ram_buffer(1956) := X"00000000";
		ram_buffer(1957) := X"00000000";
		ram_buffer(1958) := X"00000000";
		ram_buffer(1959) := X"00000000";
		ram_buffer(1960) := X"00000000";
		ram_buffer(1961) := X"00000000";
		ram_buffer(1962) := X"00000000";
		ram_buffer(1963) := X"00000000";
		ram_buffer(1964) := X"00000000";
		ram_buffer(1965) := X"00000000";
		ram_buffer(1966) := X"00000000";
		ram_buffer(1967) := X"00000000";
		ram_buffer(1968) := X"00000000";
		ram_buffer(1969) := X"00000000";
		ram_buffer(1970) := X"00000000";
		ram_buffer(1971) := X"00000000";
		ram_buffer(1972) := X"00000000";
		ram_buffer(1973) := X"00000000";
		ram_buffer(1974) := X"00000000";
		ram_buffer(1975) := X"00000000";
		ram_buffer(1976) := X"00000000";
		ram_buffer(1977) := X"00000000";
		ram_buffer(1978) := X"00000000";
		ram_buffer(1979) := X"00000000";
		ram_buffer(1980) := X"00000000";
		ram_buffer(1981) := X"00000000";
		ram_buffer(1982) := X"00000000";
		ram_buffer(1983) := X"00000000";
		ram_buffer(1984) := X"00000000";
		ram_buffer(1985) := X"00000000";
		ram_buffer(1986) := X"00000000";
		ram_buffer(1987) := X"00000000";
		ram_buffer(1988) := X"00000000";
		ram_buffer(1989) := X"00000000";
		ram_buffer(1990) := X"00000000";
		ram_buffer(1991) := X"00000000";
		ram_buffer(1992) := X"00000000";
		ram_buffer(1993) := X"00000000";
		ram_buffer(1994) := X"00000000";
		ram_buffer(1995) := X"00000000";
		ram_buffer(1996) := X"00000000";
		ram_buffer(1997) := X"00000000";
		ram_buffer(1998) := X"00000000";
		ram_buffer(1999) := X"00000000";
		ram_buffer(2000) := X"00000000";
		ram_buffer(2001) := X"00000000";
		ram_buffer(2002) := X"00000000";
		ram_buffer(2003) := X"00000000";
		ram_buffer(2004) := X"00000000";
		ram_buffer(2005) := X"00000000";
		ram_buffer(2006) := X"00000000";
		ram_buffer(2007) := X"00000000";
		ram_buffer(2008) := X"00000000";
		ram_buffer(2009) := X"00000000";
		ram_buffer(2010) := X"00000000";
		ram_buffer(2011) := X"00000000";
		ram_buffer(2012) := X"00000000";
		ram_buffer(2013) := X"00000000";
		ram_buffer(2014) := X"00000000";
		ram_buffer(2015) := X"00000000";
		ram_buffer(2016) := X"00000000";
		ram_buffer(2017) := X"00000000";
		ram_buffer(2018) := X"00000000";
		ram_buffer(2019) := X"00000000";
		ram_buffer(2020) := X"00000000";
		ram_buffer(2021) := X"00000000";
		ram_buffer(2022) := X"00000000";
		ram_buffer(2023) := X"00000000";
		ram_buffer(2024) := X"00000000";
		ram_buffer(2025) := X"00000000";
		ram_buffer(2026) := X"00000000";
		ram_buffer(2027) := X"00000000";
		ram_buffer(2028) := X"00000000";
		ram_buffer(2029) := X"00000000";
		ram_buffer(2030) := X"00000000";
		ram_buffer(2031) := X"00000000";
		ram_buffer(2032) := X"00000000";
		ram_buffer(2033) := X"00000000";
		ram_buffer(2034) := X"00000000";
		ram_buffer(2035) := X"00000000";
		ram_buffer(2036) := X"00000000";
		ram_buffer(2037) := X"00000000";
		ram_buffer(2038) := X"00000000";
		ram_buffer(2039) := X"00000000";
		ram_buffer(2040) := X"00000000";
		ram_buffer(2041) := X"00000000";
		ram_buffer(2042) := X"00000000";
		ram_buffer(2043) := X"00000000";
		ram_buffer(2044) := X"00000000";
		ram_buffer(2045) := X"00000000";
		ram_buffer(2046) := X"00000000";
		ram_buffer(2047) := X"00000000";
		ram_buffer(2048) := X"00000000";
		ram_buffer(2049) := X"00000000";
		ram_buffer(2050) := X"00000000";
		ram_buffer(2051) := X"00000000";
		ram_buffer(2052) := X"00000000";
		ram_buffer(2053) := X"00000000";
		ram_buffer(2054) := X"00000000";
		ram_buffer(2055) := X"00000000";
		ram_buffer(2056) := X"00000000";
		ram_buffer(2057) := X"00000000";
		ram_buffer(2058) := X"00000000";
		ram_buffer(2059) := X"00000000";
		ram_buffer(2060) := X"00000000";
		ram_buffer(2061) := X"00000000";
		ram_buffer(2062) := X"00000000";
		ram_buffer(2063) := X"00000000";
		ram_buffer(2064) := X"00000000";
		ram_buffer(2065) := X"00000000";
		ram_buffer(2066) := X"00000000";
		ram_buffer(2067) := X"00000000";
		ram_buffer(2068) := X"00000000";
		ram_buffer(2069) := X"00000000";
		ram_buffer(2070) := X"00000000";
		ram_buffer(2071) := X"00000000";
		ram_buffer(2072) := X"00000000";
		ram_buffer(2073) := X"00000000";
		ram_buffer(2074) := X"00000000";
		ram_buffer(2075) := X"00000000";
		ram_buffer(2076) := X"00000000";
		ram_buffer(2077) := X"00000000";
		ram_buffer(2078) := X"00000000";
		ram_buffer(2079) := X"00000000";
		ram_buffer(2080) := X"00000000";
		ram_buffer(2081) := X"00000000";
		ram_buffer(2082) := X"00000000";
		ram_buffer(2083) := X"00000000";
		ram_buffer(2084) := X"00000000";
		ram_buffer(2085) := X"00000000";
		ram_buffer(2086) := X"00000000";
		ram_buffer(2087) := X"00000000";
		ram_buffer(2088) := X"00000000";
		ram_buffer(2089) := X"00000000";
		ram_buffer(2090) := X"00000000";
		ram_buffer(2091) := X"00000000";
		ram_buffer(2092) := X"00000000";
		ram_buffer(2093) := X"00000000";
		ram_buffer(2094) := X"00000000";
		ram_buffer(2095) := X"00000000";
		ram_buffer(2096) := X"00000000";
		ram_buffer(2097) := X"00000000";
		ram_buffer(2098) := X"00000000";
		ram_buffer(2099) := X"00000000";
		ram_buffer(2100) := X"00000000";
		ram_buffer(2101) := X"00000000";
		ram_buffer(2102) := X"00000000";
		ram_buffer(2103) := X"00000000";
		ram_buffer(2104) := X"00000000";
		ram_buffer(2105) := X"00000000";
		ram_buffer(2106) := X"00000000";
		ram_buffer(2107) := X"00000000";
		ram_buffer(2108) := X"00000000";
		ram_buffer(2109) := X"00000000";
		ram_buffer(2110) := X"00000000";
		ram_buffer(2111) := X"00000000";
		ram_buffer(2112) := X"00000000";
		ram_buffer(2113) := X"00000000";
		ram_buffer(2114) := X"00000000";
		ram_buffer(2115) := X"00000000";
		ram_buffer(2116) := X"00000000";
		ram_buffer(2117) := X"00000000";
		ram_buffer(2118) := X"00000000";
		ram_buffer(2119) := X"00000000";
		ram_buffer(2120) := X"00000000";
		ram_buffer(2121) := X"00000000";
		ram_buffer(2122) := X"00000000";
		ram_buffer(2123) := X"00000000";
		ram_buffer(2124) := X"00000000";
		ram_buffer(2125) := X"00000000";
		ram_buffer(2126) := X"00000000";
		ram_buffer(2127) := X"00000000";
		ram_buffer(2128) := X"00000000";
		ram_buffer(2129) := X"00000000";
		ram_buffer(2130) := X"00000000";
		ram_buffer(2131) := X"00000000";
		ram_buffer(2132) := X"00000000";
		ram_buffer(2133) := X"00000000";
		ram_buffer(2134) := X"00000000";
		ram_buffer(2135) := X"00000000";
		ram_buffer(2136) := X"00000000";
		ram_buffer(2137) := X"00000000";
		ram_buffer(2138) := X"00000000";
		ram_buffer(2139) := X"00000000";
		ram_buffer(2140) := X"00000000";
		ram_buffer(2141) := X"00000000";
		ram_buffer(2142) := X"00000000";
		ram_buffer(2143) := X"00000000";
		ram_buffer(2144) := X"00000000";
		ram_buffer(2145) := X"00000000";
		ram_buffer(2146) := X"00000000";
		ram_buffer(2147) := X"00000000";
		ram_buffer(2148) := X"00000000";
		ram_buffer(2149) := X"00000000";
		ram_buffer(2150) := X"00000000";
		ram_buffer(2151) := X"00000000";
		ram_buffer(2152) := X"00000000";
		ram_buffer(2153) := X"00000000";
		ram_buffer(2154) := X"00000000";
		ram_buffer(2155) := X"00000000";
		ram_buffer(2156) := X"00000000";
		ram_buffer(2157) := X"00000000";
		ram_buffer(2158) := X"00000000";
		ram_buffer(2159) := X"00000000";
		ram_buffer(2160) := X"00000000";
		ram_buffer(2161) := X"00000000";
		ram_buffer(2162) := X"00000000";
		ram_buffer(2163) := X"00000000";
		ram_buffer(2164) := X"00000000";
		ram_buffer(2165) := X"00000000";
		ram_buffer(2166) := X"00000000";
		ram_buffer(2167) := X"00000000";
		ram_buffer(2168) := X"00000000";
		ram_buffer(2169) := X"00000000";
		ram_buffer(2170) := X"00000000";
		ram_buffer(2171) := X"00000000";
		ram_buffer(2172) := X"00000000";
		ram_buffer(2173) := X"00000000";
		ram_buffer(2174) := X"00000000";
		ram_buffer(2175) := X"00000000";
		ram_buffer(2176) := X"00000000";
		ram_buffer(2177) := X"00000000";
		ram_buffer(2178) := X"00000000";
		ram_buffer(2179) := X"00000000";
		ram_buffer(2180) := X"00000000";
		ram_buffer(2181) := X"00000000";
		ram_buffer(2182) := X"00000000";
		ram_buffer(2183) := X"00000000";
		ram_buffer(2184) := X"00000000";
		ram_buffer(2185) := X"00000000";
		ram_buffer(2186) := X"00000000";
		ram_buffer(2187) := X"00000000";
		ram_buffer(2188) := X"00000000";
		ram_buffer(2189) := X"00000000";
		ram_buffer(2190) := X"00000000";
		ram_buffer(2191) := X"00000000";
		ram_buffer(2192) := X"00000000";
		ram_buffer(2193) := X"00000000";
		ram_buffer(2194) := X"00000000";
		ram_buffer(2195) := X"00000000";
		ram_buffer(2196) := X"00000000";
		ram_buffer(2197) := X"00000000";
		ram_buffer(2198) := X"00000000";
		ram_buffer(2199) := X"00000000";
		ram_buffer(2200) := X"00000000";
		ram_buffer(2201) := X"00000000";
		ram_buffer(2202) := X"00000000";
		ram_buffer(2203) := X"00000000";
		ram_buffer(2204) := X"00000000";
		ram_buffer(2205) := X"00000000";
		ram_buffer(2206) := X"00000000";
		ram_buffer(2207) := X"00000000";
		ram_buffer(2208) := X"00000000";
		ram_buffer(2209) := X"00000000";
		ram_buffer(2210) := X"00000000";
		ram_buffer(2211) := X"00000000";
		ram_buffer(2212) := X"00000000";
		ram_buffer(2213) := X"00000000";
		ram_buffer(2214) := X"00000000";
		ram_buffer(2215) := X"00000000";
		ram_buffer(2216) := X"00000000";
		ram_buffer(2217) := X"00000000";
		ram_buffer(2218) := X"00000000";
		ram_buffer(2219) := X"00000000";
		ram_buffer(2220) := X"00000000";
		ram_buffer(2221) := X"00000000";
		ram_buffer(2222) := X"00000000";
		ram_buffer(2223) := X"00000000";
		ram_buffer(2224) := X"00000000";
		ram_buffer(2225) := X"00000000";
		ram_buffer(2226) := X"00000000";
		ram_buffer(2227) := X"00000000";
		ram_buffer(2228) := X"00000000";
		ram_buffer(2229) := X"00000000";
		ram_buffer(2230) := X"00000000";
		ram_buffer(2231) := X"00000000";
		ram_buffer(2232) := X"00000000";
		ram_buffer(2233) := X"00000000";
		ram_buffer(2234) := X"00000000";
		ram_buffer(2235) := X"00000000";
		ram_buffer(2236) := X"00000000";
		ram_buffer(2237) := X"00000000";
		ram_buffer(2238) := X"00000000";
		ram_buffer(2239) := X"00000000";
		ram_buffer(2240) := X"00000000";
		ram_buffer(2241) := X"00000000";
		ram_buffer(2242) := X"00000000";
		ram_buffer(2243) := X"00000000";
		ram_buffer(2244) := X"00000000";
		ram_buffer(2245) := X"00000000";
		ram_buffer(2246) := X"00000000";
		ram_buffer(2247) := X"00000000";
		ram_buffer(2248) := X"00000000";
		ram_buffer(2249) := X"00000000";
		ram_buffer(2250) := X"00000000";
		ram_buffer(2251) := X"00000000";
		ram_buffer(2252) := X"00000000";
		ram_buffer(2253) := X"00000000";
		ram_buffer(2254) := X"00000000";
		ram_buffer(2255) := X"00000000";
		ram_buffer(2256) := X"00000000";
		ram_buffer(2257) := X"00000000";
		ram_buffer(2258) := X"00000000";
		ram_buffer(2259) := X"00000000";
		ram_buffer(2260) := X"00000000";
		ram_buffer(2261) := X"00000000";
		ram_buffer(2262) := X"00000000";
		ram_buffer(2263) := X"00000000";
		ram_buffer(2264) := X"00000000";
		ram_buffer(2265) := X"00000000";
		ram_buffer(2266) := X"00000000";
		ram_buffer(2267) := X"00000000";
		ram_buffer(2268) := X"00000000";
		ram_buffer(2269) := X"00000000";
		ram_buffer(2270) := X"00000000";
		ram_buffer(2271) := X"00000000";
		ram_buffer(2272) := X"00000000";
		ram_buffer(2273) := X"00000000";
		ram_buffer(2274) := X"00000000";
		ram_buffer(2275) := X"00000000";
		ram_buffer(2276) := X"00000000";
		ram_buffer(2277) := X"00000000";
		ram_buffer(2278) := X"00000000";
		ram_buffer(2279) := X"00000000";
		ram_buffer(2280) := X"00000000";
		ram_buffer(2281) := X"00000000";
		ram_buffer(2282) := X"00000000";
		ram_buffer(2283) := X"00000000";
		ram_buffer(2284) := X"00000000";
		ram_buffer(2285) := X"00000000";
		ram_buffer(2286) := X"00000000";
		ram_buffer(2287) := X"00000000";
		ram_buffer(2288) := X"00000000";
		ram_buffer(2289) := X"00000000";
		ram_buffer(2290) := X"00000000";
		ram_buffer(2291) := X"00000000";
		ram_buffer(2292) := X"00000000";
		ram_buffer(2293) := X"00000000";
		ram_buffer(2294) := X"00000000";
		ram_buffer(2295) := X"00000000";
		ram_buffer(2296) := X"00000000";
		ram_buffer(2297) := X"00000000";
		ram_buffer(2298) := X"00000000";
		ram_buffer(2299) := X"00000000";
		ram_buffer(2300) := X"00000000";
		ram_buffer(2301) := X"00000000";
		ram_buffer(2302) := X"00000000";
		ram_buffer(2303) := X"00000000";
		ram_buffer(2304) := X"00000000";
		ram_buffer(2305) := X"00000000";
		ram_buffer(2306) := X"00000000";
		ram_buffer(2307) := X"00000000";
		ram_buffer(2308) := X"00000000";
		ram_buffer(2309) := X"00000000";
		ram_buffer(2310) := X"00000000";
		ram_buffer(2311) := X"00000000";
		ram_buffer(2312) := X"00000000";
		ram_buffer(2313) := X"00000000";
		ram_buffer(2314) := X"00000000";
		ram_buffer(2315) := X"00000000";
		ram_buffer(2316) := X"00000000";
		ram_buffer(2317) := X"00000000";
		ram_buffer(2318) := X"00000000";
		ram_buffer(2319) := X"00000000";
		ram_buffer(2320) := X"00000000";
		ram_buffer(2321) := X"00000000";
		ram_buffer(2322) := X"00000000";
		ram_buffer(2323) := X"00000000";
		ram_buffer(2324) := X"00000000";
		ram_buffer(2325) := X"00000000";
		ram_buffer(2326) := X"00000000";
		ram_buffer(2327) := X"00000000";
		ram_buffer(2328) := X"00000000";
		ram_buffer(2329) := X"00000000";
		ram_buffer(2330) := X"00000000";
		ram_buffer(2331) := X"00000000";
		ram_buffer(2332) := X"00000000";
		ram_buffer(2333) := X"00000000";
		ram_buffer(2334) := X"00000000";
		ram_buffer(2335) := X"00000000";
		ram_buffer(2336) := X"00000000";
		ram_buffer(2337) := X"00000000";
		ram_buffer(2338) := X"00000000";
		ram_buffer(2339) := X"00000000";
		ram_buffer(2340) := X"00000000";
		ram_buffer(2341) := X"00000000";
		ram_buffer(2342) := X"00000000";
		ram_buffer(2343) := X"00000000";
		ram_buffer(2344) := X"00000000";
		ram_buffer(2345) := X"00000000";
		ram_buffer(2346) := X"00000000";
		ram_buffer(2347) := X"00000000";
		ram_buffer(2348) := X"00000000";
		ram_buffer(2349) := X"00000000";
		ram_buffer(2350) := X"00000000";
		ram_buffer(2351) := X"00000000";
		ram_buffer(2352) := X"00000000";
		ram_buffer(2353) := X"00000000";
		ram_buffer(2354) := X"00000000";
		ram_buffer(2355) := X"00000000";
		ram_buffer(2356) := X"00000000";
		ram_buffer(2357) := X"00000000";
		ram_buffer(2358) := X"00000000";
		ram_buffer(2359) := X"00000000";
		ram_buffer(2360) := X"00000000";
		ram_buffer(2361) := X"00000000";
		ram_buffer(2362) := X"00000000";
		ram_buffer(2363) := X"00000000";
		ram_buffer(2364) := X"00000000";
		ram_buffer(2365) := X"00000000";
		ram_buffer(2366) := X"00000000";
		ram_buffer(2367) := X"00000000";
		ram_buffer(2368) := X"00000000";
		ram_buffer(2369) := X"00000000";
		ram_buffer(2370) := X"00000000";
		ram_buffer(2371) := X"00000000";
		ram_buffer(2372) := X"00000000";
		ram_buffer(2373) := X"00000000";
		ram_buffer(2374) := X"00000000";
		ram_buffer(2375) := X"00000000";
		ram_buffer(2376) := X"00000000";
		ram_buffer(2377) := X"00000000";
		ram_buffer(2378) := X"00000000";
		ram_buffer(2379) := X"00000000";
		ram_buffer(2380) := X"00000000";
		ram_buffer(2381) := X"00000000";
		ram_buffer(2382) := X"00000000";
		ram_buffer(2383) := X"00000000";
		ram_buffer(2384) := X"00000000";
		ram_buffer(2385) := X"00000000";
		ram_buffer(2386) := X"00000000";
		ram_buffer(2387) := X"00000000";
		ram_buffer(2388) := X"00000000";
		ram_buffer(2389) := X"00000000";
		ram_buffer(2390) := X"00000000";
		ram_buffer(2391) := X"00000000";
		ram_buffer(2392) := X"00000000";
		ram_buffer(2393) := X"00000000";
		ram_buffer(2394) := X"00000000";
		ram_buffer(2395) := X"00000000";
		ram_buffer(2396) := X"00000000";
		ram_buffer(2397) := X"00000000";
		ram_buffer(2398) := X"00000000";
		ram_buffer(2399) := X"00000000";
		ram_buffer(2400) := X"00000000";
		ram_buffer(2401) := X"00000000";
		ram_buffer(2402) := X"00000000";
		ram_buffer(2403) := X"00000000";
		ram_buffer(2404) := X"00000000";
		ram_buffer(2405) := X"00000000";
		ram_buffer(2406) := X"00000000";
		ram_buffer(2407) := X"00000000";
		ram_buffer(2408) := X"00000000";
		ram_buffer(2409) := X"00000000";
		ram_buffer(2410) := X"00000000";
		ram_buffer(2411) := X"00000000";
		ram_buffer(2412) := X"00000000";
		ram_buffer(2413) := X"00000000";
		ram_buffer(2414) := X"00000000";
		ram_buffer(2415) := X"00000000";
		ram_buffer(2416) := X"00000000";
		ram_buffer(2417) := X"00000000";
		ram_buffer(2418) := X"00000000";
		ram_buffer(2419) := X"00000000";
		ram_buffer(2420) := X"00000000";
		ram_buffer(2421) := X"00000000";
		ram_buffer(2422) := X"00000000";
		ram_buffer(2423) := X"00000000";
		ram_buffer(2424) := X"00000000";
		ram_buffer(2425) := X"00000000";
		ram_buffer(2426) := X"00000000";
		ram_buffer(2427) := X"00000000";
		ram_buffer(2428) := X"00000000";
		ram_buffer(2429) := X"00000000";
		ram_buffer(2430) := X"00000000";
		ram_buffer(2431) := X"00000000";
		ram_buffer(2432) := X"00000000";
		ram_buffer(2433) := X"00000000";
		ram_buffer(2434) := X"00000000";
		ram_buffer(2435) := X"00000000";
		ram_buffer(2436) := X"00000000";
		ram_buffer(2437) := X"00000000";
		ram_buffer(2438) := X"00000000";
		ram_buffer(2439) := X"00000000";
		ram_buffer(2440) := X"00000000";
		ram_buffer(2441) := X"00000000";
		ram_buffer(2442) := X"00000000";
		ram_buffer(2443) := X"00000000";
		ram_buffer(2444) := X"00000000";
		ram_buffer(2445) := X"00000000";
		ram_buffer(2446) := X"00000000";
		ram_buffer(2447) := X"00000000";
		ram_buffer(2448) := X"00000000";
		ram_buffer(2449) := X"00000000";
		ram_buffer(2450) := X"00000000";
		ram_buffer(2451) := X"00000000";
		ram_buffer(2452) := X"00000000";
		ram_buffer(2453) := X"00000000";
		ram_buffer(2454) := X"00000000";
		ram_buffer(2455) := X"00000000";
		ram_buffer(2456) := X"00000000";
		ram_buffer(2457) := X"00000000";
		ram_buffer(2458) := X"00000000";
		ram_buffer(2459) := X"00000000";
		ram_buffer(2460) := X"00000000";
		ram_buffer(2461) := X"00000000";
		ram_buffer(2462) := X"00000000";
		ram_buffer(2463) := X"00000000";
		ram_buffer(2464) := X"00000000";
		ram_buffer(2465) := X"00000000";
		ram_buffer(2466) := X"00000000";
		ram_buffer(2467) := X"00000000";
		ram_buffer(2468) := X"00000000";
		ram_buffer(2469) := X"00000000";
		ram_buffer(2470) := X"00000000";
		ram_buffer(2471) := X"00000000";
		ram_buffer(2472) := X"00000000";
		ram_buffer(2473) := X"00000000";
		ram_buffer(2474) := X"00000000";
		ram_buffer(2475) := X"00000000";
		ram_buffer(2476) := X"00000000";
		ram_buffer(2477) := X"00000000";
		ram_buffer(2478) := X"00000000";
		ram_buffer(2479) := X"00000000";
		ram_buffer(2480) := X"00000000";
		ram_buffer(2481) := X"00000000";
		ram_buffer(2482) := X"00000000";
		ram_buffer(2483) := X"00000000";
		ram_buffer(2484) := X"00000000";
		ram_buffer(2485) := X"00000000";
		ram_buffer(2486) := X"00000000";
		ram_buffer(2487) := X"00000000";
		ram_buffer(2488) := X"00000000";
		ram_buffer(2489) := X"00000000";
		ram_buffer(2490) := X"00000000";
		ram_buffer(2491) := X"00000000";
		ram_buffer(2492) := X"00000000";
		ram_buffer(2493) := X"00000000";
		ram_buffer(2494) := X"00000000";
		ram_buffer(2495) := X"00000000";
		ram_buffer(2496) := X"00000000";
		ram_buffer(2497) := X"00000000";
		ram_buffer(2498) := X"00000000";
		ram_buffer(2499) := X"00000000";
		ram_buffer(2500) := X"00000000";
		ram_buffer(2501) := X"00000000";
		ram_buffer(2502) := X"00000000";
		ram_buffer(2503) := X"00000000";
		ram_buffer(2504) := X"00000000";
		ram_buffer(2505) := X"00000000";
		ram_buffer(2506) := X"00000000";
		ram_buffer(2507) := X"00000000";
		ram_buffer(2508) := X"00000000";
		ram_buffer(2509) := X"00000000";
		ram_buffer(2510) := X"00000000";
		ram_buffer(2511) := X"00000000";
		ram_buffer(2512) := X"00000000";
		ram_buffer(2513) := X"00000000";
		ram_buffer(2514) := X"00000000";
		ram_buffer(2515) := X"00000000";
		ram_buffer(2516) := X"00000000";
		ram_buffer(2517) := X"00000000";
		ram_buffer(2518) := X"00000000";
		ram_buffer(2519) := X"00000000";
		ram_buffer(2520) := X"00000000";
		ram_buffer(2521) := X"00000000";
		ram_buffer(2522) := X"00000000";
		ram_buffer(2523) := X"00000000";
		ram_buffer(2524) := X"00000000";
		ram_buffer(2525) := X"00000000";
		ram_buffer(2526) := X"00000000";
		ram_buffer(2527) := X"00000000";
		ram_buffer(2528) := X"00000000";
		ram_buffer(2529) := X"00000000";
		ram_buffer(2530) := X"00000000";
		ram_buffer(2531) := X"00000000";
		ram_buffer(2532) := X"00000000";
		ram_buffer(2533) := X"00000000";
		ram_buffer(2534) := X"00000000";
		ram_buffer(2535) := X"00000000";
		ram_buffer(2536) := X"00000000";
		ram_buffer(2537) := X"00000000";
		ram_buffer(2538) := X"00000000";
		ram_buffer(2539) := X"00000000";
		ram_buffer(2540) := X"00000000";
		ram_buffer(2541) := X"00000000";
		ram_buffer(2542) := X"00000000";
		ram_buffer(2543) := X"00000000";
		ram_buffer(2544) := X"00000000";
		ram_buffer(2545) := X"00000000";
		ram_buffer(2546) := X"00000000";
		ram_buffer(2547) := X"00000000";
		ram_buffer(2548) := X"00000000";
		ram_buffer(2549) := X"00000000";
		ram_buffer(2550) := X"00000000";
		ram_buffer(2551) := X"00000000";
		ram_buffer(2552) := X"00000000";
		ram_buffer(2553) := X"00000000";
		ram_buffer(2554) := X"00000000";
		ram_buffer(2555) := X"00000000";
		ram_buffer(2556) := X"00000000";
		ram_buffer(2557) := X"00000000";
		ram_buffer(2558) := X"00000000";
		ram_buffer(2559) := X"00000000";
		ram_buffer(2560) := X"00000000";
		ram_buffer(2561) := X"00000000";
		ram_buffer(2562) := X"00000000";
		ram_buffer(2563) := X"00000000";
		ram_buffer(2564) := X"00000000";
		ram_buffer(2565) := X"00000000";
		ram_buffer(2566) := X"00000000";
		ram_buffer(2567) := X"00000000";
		ram_buffer(2568) := X"00000000";
		ram_buffer(2569) := X"00000000";
		ram_buffer(2570) := X"00000000";
		ram_buffer(2571) := X"00000000";
		ram_buffer(2572) := X"00000000";
		ram_buffer(2573) := X"00000000";
		ram_buffer(2574) := X"00000000";
		ram_buffer(2575) := X"00000000";
		ram_buffer(2576) := X"00000000";
		ram_buffer(2577) := X"00000000";
		ram_buffer(2578) := X"00000000";
		ram_buffer(2579) := X"00000000";
		ram_buffer(2580) := X"00000000";
		ram_buffer(2581) := X"00000000";
		ram_buffer(2582) := X"00000000";
		ram_buffer(2583) := X"00000000";
		ram_buffer(2584) := X"00000000";
		ram_buffer(2585) := X"00000000";
		ram_buffer(2586) := X"00000000";
		ram_buffer(2587) := X"00000000";
		ram_buffer(2588) := X"00000000";
		ram_buffer(2589) := X"00000000";
		ram_buffer(2590) := X"00000000";
		ram_buffer(2591) := X"00000000";
		ram_buffer(2592) := X"00000000";
		ram_buffer(2593) := X"00000000";
		ram_buffer(2594) := X"00000000";
		ram_buffer(2595) := X"00000000";
		ram_buffer(2596) := X"00000000";
		ram_buffer(2597) := X"00000000";
		ram_buffer(2598) := X"00000000";
		ram_buffer(2599) := X"00000000";
		ram_buffer(2600) := X"00000000";
		ram_buffer(2601) := X"00000000";
		ram_buffer(2602) := X"00000000";
		ram_buffer(2603) := X"00000000";
		ram_buffer(2604) := X"00000000";
		ram_buffer(2605) := X"00000000";
		ram_buffer(2606) := X"00000000";
		ram_buffer(2607) := X"00000000";
		ram_buffer(2608) := X"00000000";
		ram_buffer(2609) := X"00000000";
		ram_buffer(2610) := X"00000000";
		ram_buffer(2611) := X"00000000";
		ram_buffer(2612) := X"00000000";
		ram_buffer(2613) := X"00000000";
		ram_buffer(2614) := X"00000000";
		ram_buffer(2615) := X"00000000";
		ram_buffer(2616) := X"00000000";
		ram_buffer(2617) := X"00000000";
		ram_buffer(2618) := X"00000000";
		ram_buffer(2619) := X"00000000";
		ram_buffer(2620) := X"00000000";
		ram_buffer(2621) := X"00000000";
		ram_buffer(2622) := X"00000000";
		ram_buffer(2623) := X"00000000";
		ram_buffer(2624) := X"00000000";
		ram_buffer(2625) := X"00000000";
		ram_buffer(2626) := X"00000000";
		ram_buffer(2627) := X"00000000";
		ram_buffer(2628) := X"00000000";
		ram_buffer(2629) := X"00000000";
		ram_buffer(2630) := X"00000000";
		ram_buffer(2631) := X"00000000";
		ram_buffer(2632) := X"00000000";
		ram_buffer(2633) := X"00000000";
		ram_buffer(2634) := X"00000000";
		ram_buffer(2635) := X"00000000";
		ram_buffer(2636) := X"00000000";
		ram_buffer(2637) := X"00000000";
		ram_buffer(2638) := X"00000000";
		ram_buffer(2639) := X"00000000";
		ram_buffer(2640) := X"00000000";
		ram_buffer(2641) := X"00000000";
		ram_buffer(2642) := X"00000000";
		ram_buffer(2643) := X"00000000";
		ram_buffer(2644) := X"00000000";
		ram_buffer(2645) := X"00000000";
		ram_buffer(2646) := X"00000000";
		ram_buffer(2647) := X"00000000";
		ram_buffer(2648) := X"00000000";
		ram_buffer(2649) := X"00000000";
		ram_buffer(2650) := X"00000000";
		ram_buffer(2651) := X"00000000";
		ram_buffer(2652) := X"00000000";
		ram_buffer(2653) := X"00000000";
		ram_buffer(2654) := X"00000000";
		ram_buffer(2655) := X"00000000";
		ram_buffer(2656) := X"00000000";
		ram_buffer(2657) := X"00000000";
		ram_buffer(2658) := X"00000000";
		ram_buffer(2659) := X"00000000";
		ram_buffer(2660) := X"00000000";
		ram_buffer(2661) := X"00000000";
		ram_buffer(2662) := X"00000000";
		ram_buffer(2663) := X"00000000";
		ram_buffer(2664) := X"00000000";
		ram_buffer(2665) := X"00000000";
		ram_buffer(2666) := X"00000000";
		ram_buffer(2667) := X"00000000";
		ram_buffer(2668) := X"00000000";
		ram_buffer(2669) := X"00000000";
		ram_buffer(2670) := X"00000000";
		ram_buffer(2671) := X"00000000";
		ram_buffer(2672) := X"00000000";
		ram_buffer(2673) := X"00000000";
		ram_buffer(2674) := X"00000000";
		ram_buffer(2675) := X"00000000";
		ram_buffer(2676) := X"00000000";
		ram_buffer(2677) := X"00000000";
		ram_buffer(2678) := X"00000000";
		ram_buffer(2679) := X"00000000";
		ram_buffer(2680) := X"00000000";
		ram_buffer(2681) := X"00000000";
		ram_buffer(2682) := X"00000000";
		ram_buffer(2683) := X"00000000";
		ram_buffer(2684) := X"00000000";
		ram_buffer(2685) := X"00000000";
		ram_buffer(2686) := X"00000000";
		ram_buffer(2687) := X"00000000";
		ram_buffer(2688) := X"00000000";
		ram_buffer(2689) := X"00000000";
		ram_buffer(2690) := X"00000000";
		ram_buffer(2691) := X"00000000";
		ram_buffer(2692) := X"00000000";
		ram_buffer(2693) := X"00000000";
		ram_buffer(2694) := X"00000000";
		ram_buffer(2695) := X"00000000";
		ram_buffer(2696) := X"00000000";
		ram_buffer(2697) := X"00000000";
		ram_buffer(2698) := X"00000000";
		ram_buffer(2699) := X"00000000";
		ram_buffer(2700) := X"00000000";
		ram_buffer(2701) := X"00000000";
		ram_buffer(2702) := X"00000000";
		ram_buffer(2703) := X"00000000";
		ram_buffer(2704) := X"00000000";
		ram_buffer(2705) := X"00000000";
		ram_buffer(2706) := X"00000000";
		ram_buffer(2707) := X"00000000";
		ram_buffer(2708) := X"00000000";
		ram_buffer(2709) := X"00000000";
		ram_buffer(2710) := X"00000000";
		ram_buffer(2711) := X"00000000";
		ram_buffer(2712) := X"00000000";
		ram_buffer(2713) := X"00000000";
		ram_buffer(2714) := X"00000000";
		ram_buffer(2715) := X"00000000";
		ram_buffer(2716) := X"00000000";
		ram_buffer(2717) := X"00000000";
		ram_buffer(2718) := X"00000000";
		ram_buffer(2719) := X"00000000";
		ram_buffer(2720) := X"00000000";
		ram_buffer(2721) := X"00000000";
		ram_buffer(2722) := X"00000000";
		ram_buffer(2723) := X"00000000";
		ram_buffer(2724) := X"00000000";
		ram_buffer(2725) := X"00000000";
		ram_buffer(2726) := X"00000000";
		ram_buffer(2727) := X"00000000";
		ram_buffer(2728) := X"00000000";
		ram_buffer(2729) := X"00000000";
		ram_buffer(2730) := X"00000000";
		ram_buffer(2731) := X"00000000";
		ram_buffer(2732) := X"00000000";
		ram_buffer(2733) := X"00000000";
		ram_buffer(2734) := X"00000000";
		ram_buffer(2735) := X"00000000";
		ram_buffer(2736) := X"00000000";
		ram_buffer(2737) := X"00000000";
		ram_buffer(2738) := X"00000000";
		ram_buffer(2739) := X"00000000";
		ram_buffer(2740) := X"00000000";
		ram_buffer(2741) := X"00000000";
		ram_buffer(2742) := X"00000000";
		ram_buffer(2743) := X"00000000";
		ram_buffer(2744) := X"00000000";
		ram_buffer(2745) := X"00000000";
		ram_buffer(2746) := X"00000000";
		ram_buffer(2747) := X"00000000";
		ram_buffer(2748) := X"00000000";
		ram_buffer(2749) := X"00000000";
		ram_buffer(2750) := X"00000000";
		ram_buffer(2751) := X"00000000";
		ram_buffer(2752) := X"00000000";
		ram_buffer(2753) := X"00000000";
		ram_buffer(2754) := X"00000000";
		ram_buffer(2755) := X"00000000";
		ram_buffer(2756) := X"00000000";
		ram_buffer(2757) := X"00000000";
		ram_buffer(2758) := X"00000000";
		ram_buffer(2759) := X"00000000";
		ram_buffer(2760) := X"00000000";
		ram_buffer(2761) := X"00000000";
		ram_buffer(2762) := X"00000000";
		ram_buffer(2763) := X"00000000";
		ram_buffer(2764) := X"00000000";
		ram_buffer(2765) := X"00000000";
		ram_buffer(2766) := X"00000000";
		ram_buffer(2767) := X"00000000";
		ram_buffer(2768) := X"00000000";
		ram_buffer(2769) := X"00000000";
		ram_buffer(2770) := X"00000000";
		ram_buffer(2771) := X"00000000";
		ram_buffer(2772) := X"00000000";
		ram_buffer(2773) := X"00000000";
		ram_buffer(2774) := X"00000000";
		ram_buffer(2775) := X"00000000";
		ram_buffer(2776) := X"00000000";
		ram_buffer(2777) := X"00000000";
		ram_buffer(2778) := X"00000000";
		ram_buffer(2779) := X"00000000";
		ram_buffer(2780) := X"00000000";
		ram_buffer(2781) := X"00000000";
		ram_buffer(2782) := X"00000000";
		ram_buffer(2783) := X"00000000";
		ram_buffer(2784) := X"00000000";
		ram_buffer(2785) := X"00000000";
		ram_buffer(2786) := X"00000000";
		ram_buffer(2787) := X"00000000";
		ram_buffer(2788) := X"00000000";
		ram_buffer(2789) := X"00000000";
		ram_buffer(2790) := X"00000000";
		ram_buffer(2791) := X"00000000";
		ram_buffer(2792) := X"00000000";
		ram_buffer(2793) := X"00000000";
		ram_buffer(2794) := X"00000000";
		ram_buffer(2795) := X"00000000";
		ram_buffer(2796) := X"00000000";
		ram_buffer(2797) := X"00000000";
		ram_buffer(2798) := X"00000000";
		ram_buffer(2799) := X"00000000";
		ram_buffer(2800) := X"00000000";
		ram_buffer(2801) := X"00000000";
		ram_buffer(2802) := X"00000000";
		ram_buffer(2803) := X"00000000";
		ram_buffer(2804) := X"00000000";
		ram_buffer(2805) := X"00000000";
		ram_buffer(2806) := X"00000000";
		ram_buffer(2807) := X"00000000";
		ram_buffer(2808) := X"00000000";
		ram_buffer(2809) := X"00000000";
		ram_buffer(2810) := X"00000000";
		ram_buffer(2811) := X"00000000";
		ram_buffer(2812) := X"00000000";
		ram_buffer(2813) := X"00000000";
		ram_buffer(2814) := X"00000000";
		ram_buffer(2815) := X"00000000";
		ram_buffer(2816) := X"00000000";
		ram_buffer(2817) := X"00000000";
		ram_buffer(2818) := X"00000000";
		ram_buffer(2819) := X"00000000";
		ram_buffer(2820) := X"00000000";
		ram_buffer(2821) := X"00000000";
		ram_buffer(2822) := X"00000000";
		ram_buffer(2823) := X"00000000";
		ram_buffer(2824) := X"00000000";
		ram_buffer(2825) := X"00000000";
		ram_buffer(2826) := X"00000000";
		ram_buffer(2827) := X"00000000";
		ram_buffer(2828) := X"00000000";
		ram_buffer(2829) := X"00000000";
		ram_buffer(2830) := X"00000000";
		ram_buffer(2831) := X"00000000";
		ram_buffer(2832) := X"00000000";
		ram_buffer(2833) := X"00000000";
		ram_buffer(2834) := X"00000000";
		ram_buffer(2835) := X"00000000";
		ram_buffer(2836) := X"00000000";
		ram_buffer(2837) := X"00000000";
		ram_buffer(2838) := X"00000000";
		ram_buffer(2839) := X"00000000";
		ram_buffer(2840) := X"00000000";
		ram_buffer(2841) := X"00000000";
		ram_buffer(2842) := X"00000000";
		ram_buffer(2843) := X"00000000";
		ram_buffer(2844) := X"00000000";
		ram_buffer(2845) := X"00000000";
		ram_buffer(2846) := X"00000000";
		ram_buffer(2847) := X"00000000";
		ram_buffer(2848) := X"00000000";
		ram_buffer(2849) := X"00000000";
		ram_buffer(2850) := X"00000000";
		ram_buffer(2851) := X"00000000";
		ram_buffer(2852) := X"00000000";
		ram_buffer(2853) := X"00000000";
		ram_buffer(2854) := X"00000000";
		ram_buffer(2855) := X"00000000";
		ram_buffer(2856) := X"00000000";
		ram_buffer(2857) := X"00000000";
		ram_buffer(2858) := X"00000000";
		ram_buffer(2859) := X"00000000";
		ram_buffer(2860) := X"00000000";
		ram_buffer(2861) := X"00000000";
		ram_buffer(2862) := X"00000000";
		ram_buffer(2863) := X"00000000";
		ram_buffer(2864) := X"00000000";
		ram_buffer(2865) := X"00000000";
		ram_buffer(2866) := X"00000000";
		ram_buffer(2867) := X"00000000";
		ram_buffer(2868) := X"00000000";
		ram_buffer(2869) := X"00000000";
		ram_buffer(2870) := X"00000000";
		ram_buffer(2871) := X"00000000";
		ram_buffer(2872) := X"00000000";
		ram_buffer(2873) := X"00000000";
		ram_buffer(2874) := X"00000000";
		ram_buffer(2875) := X"00000000";
		ram_buffer(2876) := X"00000000";
		ram_buffer(2877) := X"00000000";
		ram_buffer(2878) := X"00000000";
		ram_buffer(2879) := X"00000000";
		ram_buffer(2880) := X"00000000";
		ram_buffer(2881) := X"00000000";
		ram_buffer(2882) := X"00000000";
		ram_buffer(2883) := X"00000000";
		ram_buffer(2884) := X"00000000";
		ram_buffer(2885) := X"00000000";
		ram_buffer(2886) := X"00000000";
		ram_buffer(2887) := X"00000000";
		ram_buffer(2888) := X"00000000";
		ram_buffer(2889) := X"00000000";
		ram_buffer(2890) := X"00000000";
		ram_buffer(2891) := X"00000000";
		ram_buffer(2892) := X"00000000";
		ram_buffer(2893) := X"00000000";
		ram_buffer(2894) := X"00000000";
		ram_buffer(2895) := X"00000000";
		ram_buffer(2896) := X"00000000";
		ram_buffer(2897) := X"00000000";
		ram_buffer(2898) := X"00000000";
		ram_buffer(2899) := X"00000000";
		ram_buffer(2900) := X"00000000";
		ram_buffer(2901) := X"00000000";
		ram_buffer(2902) := X"00000000";
		ram_buffer(2903) := X"00000000";
		ram_buffer(2904) := X"00000000";
		ram_buffer(2905) := X"00000000";
		ram_buffer(2906) := X"00000000";
		ram_buffer(2907) := X"00000000";
		ram_buffer(2908) := X"00000000";
		ram_buffer(2909) := X"00000000";
		ram_buffer(2910) := X"00000000";
		ram_buffer(2911) := X"00000000";
		ram_buffer(2912) := X"00000000";
		ram_buffer(2913) := X"00000000";
		ram_buffer(2914) := X"00000000";
		ram_buffer(2915) := X"00000000";
		ram_buffer(2916) := X"00000000";
		ram_buffer(2917) := X"00000000";
		ram_buffer(2918) := X"00000000";
		ram_buffer(2919) := X"00000000";
		ram_buffer(2920) := X"00000000";
		ram_buffer(2921) := X"00000000";
		ram_buffer(2922) := X"00000000";
		ram_buffer(2923) := X"00000000";
		ram_buffer(2924) := X"00000000";
		ram_buffer(2925) := X"00000000";
		ram_buffer(2926) := X"00000000";
		ram_buffer(2927) := X"00000000";
		ram_buffer(2928) := X"00000000";
		ram_buffer(2929) := X"00000000";
		ram_buffer(2930) := X"00000000";
		ram_buffer(2931) := X"00000000";
		ram_buffer(2932) := X"00000000";
		ram_buffer(2933) := X"00000000";
		ram_buffer(2934) := X"00000000";
		ram_buffer(2935) := X"00000000";
		ram_buffer(2936) := X"00000000";
		ram_buffer(2937) := X"00000000";
		ram_buffer(2938) := X"00000000";
		ram_buffer(2939) := X"00000000";
		ram_buffer(2940) := X"00000000";
		ram_buffer(2941) := X"00000000";
		ram_buffer(2942) := X"00000000";
		ram_buffer(2943) := X"00000000";
		ram_buffer(2944) := X"00000000";
		ram_buffer(2945) := X"00000000";
		ram_buffer(2946) := X"00000000";
		ram_buffer(2947) := X"00000000";
		ram_buffer(2948) := X"00000000";
		ram_buffer(2949) := X"00000000";
		ram_buffer(2950) := X"00000000";
		ram_buffer(2951) := X"00000000";
		ram_buffer(2952) := X"00000000";
		ram_buffer(2953) := X"00000000";
		ram_buffer(2954) := X"00000000";
		ram_buffer(2955) := X"00000000";
		ram_buffer(2956) := X"00000000";
		ram_buffer(2957) := X"00000000";
		ram_buffer(2958) := X"00000000";
		ram_buffer(2959) := X"00000000";
		ram_buffer(2960) := X"00000000";
		ram_buffer(2961) := X"00000000";
		ram_buffer(2962) := X"00000000";
		ram_buffer(2963) := X"00000000";
		ram_buffer(2964) := X"00000000";
		ram_buffer(2965) := X"00000000";
		ram_buffer(2966) := X"00000000";
		ram_buffer(2967) := X"00000000";
		ram_buffer(2968) := X"00000000";
		ram_buffer(2969) := X"00000000";
		ram_buffer(2970) := X"00000000";
		ram_buffer(2971) := X"00000000";
		ram_buffer(2972) := X"00000000";
		ram_buffer(2973) := X"00000000";
		ram_buffer(2974) := X"00000000";
		ram_buffer(2975) := X"00000000";
		ram_buffer(2976) := X"00000000";
		ram_buffer(2977) := X"00000000";
		ram_buffer(2978) := X"00000000";
		ram_buffer(2979) := X"00000000";
		ram_buffer(2980) := X"00000000";
		ram_buffer(2981) := X"00000000";
		ram_buffer(2982) := X"00000000";
		ram_buffer(2983) := X"00000000";
		ram_buffer(2984) := X"00000000";
		ram_buffer(2985) := X"00000000";
		ram_buffer(2986) := X"00000000";
		ram_buffer(2987) := X"00000000";
		ram_buffer(2988) := X"00000000";
		ram_buffer(2989) := X"00000000";
		ram_buffer(2990) := X"00000000";
		ram_buffer(2991) := X"00000000";
		ram_buffer(2992) := X"00000000";
		ram_buffer(2993) := X"00000000";
		ram_buffer(2994) := X"00000000";
		ram_buffer(2995) := X"00000000";
		ram_buffer(2996) := X"00000000";
		ram_buffer(2997) := X"00000000";
		ram_buffer(2998) := X"00000000";
		ram_buffer(2999) := X"00000000";
		ram_buffer(3000) := X"00000000";
		ram_buffer(3001) := X"00000000";
		ram_buffer(3002) := X"00000000";
		ram_buffer(3003) := X"00000000";
		ram_buffer(3004) := X"00000000";
		ram_buffer(3005) := X"00000000";
		ram_buffer(3006) := X"00000000";
		ram_buffer(3007) := X"00000000";
		ram_buffer(3008) := X"00000000";
		ram_buffer(3009) := X"00000000";
		ram_buffer(3010) := X"00000000";
		ram_buffer(3011) := X"00000000";
		ram_buffer(3012) := X"00000000";
		ram_buffer(3013) := X"00000000";
		ram_buffer(3014) := X"00000000";
		ram_buffer(3015) := X"00000000";
		ram_buffer(3016) := X"00000000";
		ram_buffer(3017) := X"00000000";
		ram_buffer(3018) := X"00000000";
		ram_buffer(3019) := X"00000000";
		ram_buffer(3020) := X"00000000";
		ram_buffer(3021) := X"00000000";
		ram_buffer(3022) := X"00000000";
		ram_buffer(3023) := X"00000000";
		ram_buffer(3024) := X"00000000";
		ram_buffer(3025) := X"00000000";
		ram_buffer(3026) := X"00000000";
		ram_buffer(3027) := X"00000000";
		ram_buffer(3028) := X"00000000";
		ram_buffer(3029) := X"00000000";
		ram_buffer(3030) := X"00000000";
		ram_buffer(3031) := X"00000000";
		ram_buffer(3032) := X"00000000";
		ram_buffer(3033) := X"00000000";
		ram_buffer(3034) := X"00000000";
		ram_buffer(3035) := X"00000000";
		ram_buffer(3036) := X"00000000";
		ram_buffer(3037) := X"00000000";
		ram_buffer(3038) := X"00000000";
		ram_buffer(3039) := X"00000000";
		ram_buffer(3040) := X"00000000";
		ram_buffer(3041) := X"00000000";
		ram_buffer(3042) := X"00000000";
		ram_buffer(3043) := X"00000000";
		ram_buffer(3044) := X"00000000";
		ram_buffer(3045) := X"00000000";
		ram_buffer(3046) := X"00000000";
		ram_buffer(3047) := X"00000000";
		ram_buffer(3048) := X"00000000";
		ram_buffer(3049) := X"00000000";
		ram_buffer(3050) := X"00000000";
		ram_buffer(3051) := X"00000000";
		ram_buffer(3052) := X"00000000";
		ram_buffer(3053) := X"00000000";
		ram_buffer(3054) := X"00000000";
		ram_buffer(3055) := X"00000000";
		ram_buffer(3056) := X"00000000";
		ram_buffer(3057) := X"00000000";
		ram_buffer(3058) := X"00000000";
		ram_buffer(3059) := X"00000000";
		ram_buffer(3060) := X"00000000";
		ram_buffer(3061) := X"00000000";
		ram_buffer(3062) := X"00000000";
		ram_buffer(3063) := X"00000000";
		ram_buffer(3064) := X"00000000";
		ram_buffer(3065) := X"00000000";
		ram_buffer(3066) := X"00000000";
		ram_buffer(3067) := X"00000000";
		ram_buffer(3068) := X"00000000";
		ram_buffer(3069) := X"00000000";
		ram_buffer(3070) := X"00000000";
		ram_buffer(3071) := X"00000000";
		ram_buffer(3072) := X"00000000";
		ram_buffer(3073) := X"00000000";
		ram_buffer(3074) := X"00000000";
		ram_buffer(3075) := X"00000000";
		ram_buffer(3076) := X"00000000";
		ram_buffer(3077) := X"00000000";
		ram_buffer(3078) := X"00000000";
		ram_buffer(3079) := X"00000000";
		ram_buffer(3080) := X"00000000";
		ram_buffer(3081) := X"00000000";
		ram_buffer(3082) := X"00000000";
		ram_buffer(3083) := X"00000000";
		ram_buffer(3084) := X"00000000";
		ram_buffer(3085) := X"00000000";
		ram_buffer(3086) := X"00000000";
		ram_buffer(3087) := X"00000000";
		ram_buffer(3088) := X"00000000";
		ram_buffer(3089) := X"00000000";
		ram_buffer(3090) := X"00000000";
		ram_buffer(3091) := X"00000000";
		ram_buffer(3092) := X"00000000";
		ram_buffer(3093) := X"00000000";
		ram_buffer(3094) := X"00000000";
		ram_buffer(3095) := X"00000000";
		ram_buffer(3096) := X"00000000";
		ram_buffer(3097) := X"00000000";
		ram_buffer(3098) := X"00000000";
		ram_buffer(3099) := X"00000000";
		ram_buffer(3100) := X"00000000";
		ram_buffer(3101) := X"00000000";
		ram_buffer(3102) := X"00000000";
		ram_buffer(3103) := X"00000000";
		ram_buffer(3104) := X"00000000";
		ram_buffer(3105) := X"00000000";
		ram_buffer(3106) := X"00000000";
		ram_buffer(3107) := X"00000000";
		ram_buffer(3108) := X"00000000";
		ram_buffer(3109) := X"00000000";
		ram_buffer(3110) := X"00000000";
		ram_buffer(3111) := X"00000000";
		ram_buffer(3112) := X"00000000";
		ram_buffer(3113) := X"00000000";
		ram_buffer(3114) := X"00000000";
		ram_buffer(3115) := X"00000000";
		ram_buffer(3116) := X"00000000";
		ram_buffer(3117) := X"00000000";
		ram_buffer(3118) := X"00000000";
		ram_buffer(3119) := X"00000000";
		ram_buffer(3120) := X"00000000";
		ram_buffer(3121) := X"00000000";
		ram_buffer(3122) := X"00000000";
		ram_buffer(3123) := X"00000000";
		ram_buffer(3124) := X"00000000";
		ram_buffer(3125) := X"00000000";
		ram_buffer(3126) := X"00000000";
		ram_buffer(3127) := X"00000000";
		ram_buffer(3128) := X"00000000";
		ram_buffer(3129) := X"00000000";
		ram_buffer(3130) := X"00000000";
		ram_buffer(3131) := X"00000000";
		ram_buffer(3132) := X"00000000";
		ram_buffer(3133) := X"00000000";
		ram_buffer(3134) := X"00000000";
		ram_buffer(3135) := X"00000000";
		ram_buffer(3136) := X"00000000";
		ram_buffer(3137) := X"00000000";
		ram_buffer(3138) := X"00000000";
		ram_buffer(3139) := X"00000000";
		ram_buffer(3140) := X"00000000";
		ram_buffer(3141) := X"00000000";
		ram_buffer(3142) := X"00000000";
		ram_buffer(3143) := X"00000000";
		ram_buffer(3144) := X"00000000";
		ram_buffer(3145) := X"00000000";
		ram_buffer(3146) := X"00000000";
		ram_buffer(3147) := X"00000000";
		ram_buffer(3148) := X"00000000";
		ram_buffer(3149) := X"00000000";
		ram_buffer(3150) := X"00000000";
		ram_buffer(3151) := X"00000000";
		ram_buffer(3152) := X"00000000";
		ram_buffer(3153) := X"00000000";
		ram_buffer(3154) := X"00000000";
		ram_buffer(3155) := X"00000000";
		ram_buffer(3156) := X"00000000";
		ram_buffer(3157) := X"00000000";
		ram_buffer(3158) := X"00000000";
		ram_buffer(3159) := X"00000000";
		ram_buffer(3160) := X"00000000";
		ram_buffer(3161) := X"00000000";
		ram_buffer(3162) := X"00000000";
		ram_buffer(3163) := X"00000000";
		ram_buffer(3164) := X"00000000";
		ram_buffer(3165) := X"00000000";
		ram_buffer(3166) := X"00000000";
		ram_buffer(3167) := X"00000000";
		ram_buffer(3168) := X"00000000";
		ram_buffer(3169) := X"00000000";
		ram_buffer(3170) := X"00000000";
		ram_buffer(3171) := X"00000000";
		ram_buffer(3172) := X"00000000";
		ram_buffer(3173) := X"00000000";
		ram_buffer(3174) := X"00000000";
		ram_buffer(3175) := X"00000000";
		ram_buffer(3176) := X"00000000";
		ram_buffer(3177) := X"00000000";
		ram_buffer(3178) := X"00000000";
		ram_buffer(3179) := X"00000000";
		ram_buffer(3180) := X"00000000";
		ram_buffer(3181) := X"00000000";
		ram_buffer(3182) := X"00000000";
		ram_buffer(3183) := X"00000000";
		ram_buffer(3184) := X"00000000";
		ram_buffer(3185) := X"00000000";
		ram_buffer(3186) := X"00000000";
		ram_buffer(3187) := X"00000000";
		ram_buffer(3188) := X"00000000";
		ram_buffer(3189) := X"00000000";
		ram_buffer(3190) := X"00000000";
		ram_buffer(3191) := X"00000000";
		ram_buffer(3192) := X"00000000";
		ram_buffer(3193) := X"00000000";
		ram_buffer(3194) := X"00000000";
		ram_buffer(3195) := X"00000000";
		ram_buffer(3196) := X"00000000";
		ram_buffer(3197) := X"00000000";
		ram_buffer(3198) := X"00000000";
		ram_buffer(3199) := X"00000000";
		ram_buffer(3200) := X"00000000";
		ram_buffer(3201) := X"00000000";
		ram_buffer(3202) := X"00000000";
		ram_buffer(3203) := X"00000000";
		ram_buffer(3204) := X"00000000";
		ram_buffer(3205) := X"00000000";
		ram_buffer(3206) := X"00000000";
		ram_buffer(3207) := X"00000000";
		ram_buffer(3208) := X"00000000";
		ram_buffer(3209) := X"00000000";
		ram_buffer(3210) := X"00000000";
		ram_buffer(3211) := X"00000000";
		ram_buffer(3212) := X"00000000";
		ram_buffer(3213) := X"00000000";
		ram_buffer(3214) := X"00000000";
		ram_buffer(3215) := X"00000000";
		ram_buffer(3216) := X"00000000";
		ram_buffer(3217) := X"00000000";
		ram_buffer(3218) := X"00000000";
		ram_buffer(3219) := X"00000000";
		ram_buffer(3220) := X"00000000";
		ram_buffer(3221) := X"00000000";
		ram_buffer(3222) := X"00000000";
		ram_buffer(3223) := X"00000000";
		ram_buffer(3224) := X"00000000";
		ram_buffer(3225) := X"00000000";
		ram_buffer(3226) := X"00000000";
		ram_buffer(3227) := X"00000000";
		ram_buffer(3228) := X"00000000";
		ram_buffer(3229) := X"00000000";
		ram_buffer(3230) := X"00000000";
		ram_buffer(3231) := X"00000000";
		ram_buffer(3232) := X"00000000";
		ram_buffer(3233) := X"00000000";
		ram_buffer(3234) := X"00000000";
		ram_buffer(3235) := X"00000000";
		ram_buffer(3236) := X"00000000";
		ram_buffer(3237) := X"00000000";
		ram_buffer(3238) := X"00000000";
		ram_buffer(3239) := X"00000000";
		ram_buffer(3240) := X"00000000";
		ram_buffer(3241) := X"00000000";
		ram_buffer(3242) := X"00000000";
		ram_buffer(3243) := X"00000000";
		ram_buffer(3244) := X"00000000";
		ram_buffer(3245) := X"00000000";
		ram_buffer(3246) := X"00000000";
		ram_buffer(3247) := X"00000000";
		ram_buffer(3248) := X"00000000";
		ram_buffer(3249) := X"00000000";
		ram_buffer(3250) := X"00000000";
		ram_buffer(3251) := X"00000000";
		ram_buffer(3252) := X"00000000";
		ram_buffer(3253) := X"00000000";
		ram_buffer(3254) := X"00000000";
		ram_buffer(3255) := X"00000000";
		ram_buffer(3256) := X"00000000";
		ram_buffer(3257) := X"00000000";
		ram_buffer(3258) := X"00000000";
		ram_buffer(3259) := X"00000000";
		ram_buffer(3260) := X"00000000";
		ram_buffer(3261) := X"00000000";
		ram_buffer(3262) := X"00000000";
		ram_buffer(3263) := X"00000000";
		ram_buffer(3264) := X"00000000";
		ram_buffer(3265) := X"00000000";
		ram_buffer(3266) := X"00000000";
		ram_buffer(3267) := X"00000000";
		ram_buffer(3268) := X"00000000";
		ram_buffer(3269) := X"00000000";
		ram_buffer(3270) := X"00000000";
		ram_buffer(3271) := X"00000000";
		ram_buffer(3272) := X"00000000";
		ram_buffer(3273) := X"00000000";
		ram_buffer(3274) := X"00000000";
		ram_buffer(3275) := X"00000000";
		ram_buffer(3276) := X"00000000";
		ram_buffer(3277) := X"00000000";
		ram_buffer(3278) := X"00000000";
		ram_buffer(3279) := X"00000000";
		ram_buffer(3280) := X"00000000";
		ram_buffer(3281) := X"00000000";
		ram_buffer(3282) := X"00000000";
		ram_buffer(3283) := X"00000000";
		ram_buffer(3284) := X"00000000";
		ram_buffer(3285) := X"00000000";
		ram_buffer(3286) := X"00000000";
		ram_buffer(3287) := X"00000000";
		ram_buffer(3288) := X"00000000";
		ram_buffer(3289) := X"00000000";
		ram_buffer(3290) := X"00000000";
		ram_buffer(3291) := X"00000000";
		ram_buffer(3292) := X"00000000";
		ram_buffer(3293) := X"00000000";
		ram_buffer(3294) := X"00000000";
		ram_buffer(3295) := X"00000000";
		ram_buffer(3296) := X"00000000";
		ram_buffer(3297) := X"00000000";
		ram_buffer(3298) := X"00000000";
		ram_buffer(3299) := X"00000000";
		ram_buffer(3300) := X"00000000";
		ram_buffer(3301) := X"00000000";
		ram_buffer(3302) := X"00000000";
		ram_buffer(3303) := X"00000000";
		ram_buffer(3304) := X"00000000";
		ram_buffer(3305) := X"00000000";
		ram_buffer(3306) := X"00000000";
		ram_buffer(3307) := X"00000000";
		ram_buffer(3308) := X"00000000";
		ram_buffer(3309) := X"00000000";
		ram_buffer(3310) := X"00000000";
		ram_buffer(3311) := X"00000000";
		ram_buffer(3312) := X"00000000";
		ram_buffer(3313) := X"00000000";
		ram_buffer(3314) := X"00000000";
		ram_buffer(3315) := X"00000000";
		ram_buffer(3316) := X"00000000";
		ram_buffer(3317) := X"00000000";
		ram_buffer(3318) := X"00000000";
		ram_buffer(3319) := X"00000000";
		ram_buffer(3320) := X"00000000";
		ram_buffer(3321) := X"00000000";
		ram_buffer(3322) := X"00000000";
		ram_buffer(3323) := X"00000000";
		ram_buffer(3324) := X"00000000";
		ram_buffer(3325) := X"00000000";
		ram_buffer(3326) := X"00000000";
		ram_buffer(3327) := X"00000000";
		ram_buffer(3328) := X"00000000";
		ram_buffer(3329) := X"00000000";
		ram_buffer(3330) := X"00000000";
		ram_buffer(3331) := X"00000000";
		ram_buffer(3332) := X"00000000";
		ram_buffer(3333) := X"00000000";
		ram_buffer(3334) := X"00000000";
		ram_buffer(3335) := X"00000000";
		ram_buffer(3336) := X"00000000";
		ram_buffer(3337) := X"00000000";
		ram_buffer(3338) := X"00000000";
		ram_buffer(3339) := X"00000000";
		ram_buffer(3340) := X"00000000";
		ram_buffer(3341) := X"00000000";
		ram_buffer(3342) := X"00000000";
		ram_buffer(3343) := X"00000000";
		ram_buffer(3344) := X"00000000";
		ram_buffer(3345) := X"00000000";
		ram_buffer(3346) := X"00000000";
		ram_buffer(3347) := X"00000000";
		ram_buffer(3348) := X"00000000";
		ram_buffer(3349) := X"00000000";
		ram_buffer(3350) := X"00000000";
		ram_buffer(3351) := X"00000000";
		ram_buffer(3352) := X"00000000";
		ram_buffer(3353) := X"00000000";
		ram_buffer(3354) := X"00000000";
		ram_buffer(3355) := X"00000000";
		ram_buffer(3356) := X"00000000";
		ram_buffer(3357) := X"00000000";
		ram_buffer(3358) := X"00000000";
		ram_buffer(3359) := X"00000000";
		ram_buffer(3360) := X"00000000";
		ram_buffer(3361) := X"00000000";
		ram_buffer(3362) := X"00000000";
		ram_buffer(3363) := X"00000000";
		ram_buffer(3364) := X"00000000";
		ram_buffer(3365) := X"00000000";
		ram_buffer(3366) := X"00000000";
		ram_buffer(3367) := X"00000000";
		ram_buffer(3368) := X"00000000";
		ram_buffer(3369) := X"00000000";
		ram_buffer(3370) := X"00000000";
		ram_buffer(3371) := X"00000000";
		ram_buffer(3372) := X"00000000";
		ram_buffer(3373) := X"00000000";
		ram_buffer(3374) := X"00000000";
		ram_buffer(3375) := X"00000000";
		ram_buffer(3376) := X"00000000";
		ram_buffer(3377) := X"00000000";
		ram_buffer(3378) := X"00000000";
		ram_buffer(3379) := X"00000000";
		ram_buffer(3380) := X"00000000";
		ram_buffer(3381) := X"00000000";
		ram_buffer(3382) := X"00000000";
		ram_buffer(3383) := X"00000000";
		ram_buffer(3384) := X"00000000";
		ram_buffer(3385) := X"00000000";
		ram_buffer(3386) := X"00000000";
		ram_buffer(3387) := X"00000000";
		ram_buffer(3388) := X"00000000";
		ram_buffer(3389) := X"00000000";
		ram_buffer(3390) := X"00000000";
		ram_buffer(3391) := X"00000000";
		ram_buffer(3392) := X"00000000";
		ram_buffer(3393) := X"00000000";
		ram_buffer(3394) := X"00000000";
		ram_buffer(3395) := X"00000000";
		ram_buffer(3396) := X"00000000";
		ram_buffer(3397) := X"00000000";
		ram_buffer(3398) := X"00000000";
		ram_buffer(3399) := X"00000000";
		ram_buffer(3400) := X"00000000";
		ram_buffer(3401) := X"00000000";
		ram_buffer(3402) := X"00000000";
		ram_buffer(3403) := X"00000000";
		ram_buffer(3404) := X"00000000";
		ram_buffer(3405) := X"00000000";
		ram_buffer(3406) := X"00000000";
		ram_buffer(3407) := X"00000000";
		ram_buffer(3408) := X"00000000";
		ram_buffer(3409) := X"00000000";
		ram_buffer(3410) := X"00000000";
		ram_buffer(3411) := X"00000000";
		ram_buffer(3412) := X"00000000";
		ram_buffer(3413) := X"00000000";
		ram_buffer(3414) := X"00000000";
		ram_buffer(3415) := X"00000000";
		ram_buffer(3416) := X"00000000";
		ram_buffer(3417) := X"00000000";
		ram_buffer(3418) := X"00000000";
		ram_buffer(3419) := X"00000000";
		ram_buffer(3420) := X"00000000";
		ram_buffer(3421) := X"00000000";
		ram_buffer(3422) := X"00000000";
		ram_buffer(3423) := X"00000000";
		ram_buffer(3424) := X"00000000";
		ram_buffer(3425) := X"00000000";
		ram_buffer(3426) := X"00000000";
		ram_buffer(3427) := X"00000000";
		ram_buffer(3428) := X"00000000";
		ram_buffer(3429) := X"00000000";
		ram_buffer(3430) := X"00000000";
		ram_buffer(3431) := X"00000000";
		ram_buffer(3432) := X"00000000";
		ram_buffer(3433) := X"00000000";
		ram_buffer(3434) := X"00000000";
		ram_buffer(3435) := X"00000000";
		ram_buffer(3436) := X"00000000";
		ram_buffer(3437) := X"00000000";
		ram_buffer(3438) := X"00000000";
		ram_buffer(3439) := X"00000000";
		ram_buffer(3440) := X"00000000";
		ram_buffer(3441) := X"00000000";
		ram_buffer(3442) := X"00000000";
		ram_buffer(3443) := X"00000000";
		ram_buffer(3444) := X"00000000";
		ram_buffer(3445) := X"00000000";
		ram_buffer(3446) := X"00000000";
		ram_buffer(3447) := X"00000000";
		ram_buffer(3448) := X"00000000";
		ram_buffer(3449) := X"00000000";
		ram_buffer(3450) := X"00000000";
		ram_buffer(3451) := X"00000000";
		ram_buffer(3452) := X"00000000";
		ram_buffer(3453) := X"00000000";
		ram_buffer(3454) := X"00000000";
		ram_buffer(3455) := X"00000000";
		ram_buffer(3456) := X"00000000";
		ram_buffer(3457) := X"00000000";
		ram_buffer(3458) := X"00000000";
		ram_buffer(3459) := X"00000000";
		ram_buffer(3460) := X"00000000";
		ram_buffer(3461) := X"00000000";
		ram_buffer(3462) := X"00000000";
		ram_buffer(3463) := X"00000000";
		ram_buffer(3464) := X"00000000";
		ram_buffer(3465) := X"00000000";
		ram_buffer(3466) := X"00000000";
		ram_buffer(3467) := X"00000000";
		ram_buffer(3468) := X"00000000";
		ram_buffer(3469) := X"00000000";
		ram_buffer(3470) := X"00000000";
		ram_buffer(3471) := X"00000000";
		ram_buffer(3472) := X"00000000";
		ram_buffer(3473) := X"00000000";
		ram_buffer(3474) := X"00000000";
		ram_buffer(3475) := X"00000000";
		ram_buffer(3476) := X"00000000";
		ram_buffer(3477) := X"00000000";
		ram_buffer(3478) := X"00000000";
		ram_buffer(3479) := X"00000000";
		ram_buffer(3480) := X"00000000";
		ram_buffer(3481) := X"00000000";
		ram_buffer(3482) := X"00000000";
		ram_buffer(3483) := X"00000000";
		ram_buffer(3484) := X"00000000";
		ram_buffer(3485) := X"00000000";
		ram_buffer(3486) := X"00000000";
		ram_buffer(3487) := X"00000000";
		ram_buffer(3488) := X"00000000";
		ram_buffer(3489) := X"00000000";
		ram_buffer(3490) := X"00000000";
		ram_buffer(3491) := X"00000000";
		ram_buffer(3492) := X"00000000";
		ram_buffer(3493) := X"00000000";
		ram_buffer(3494) := X"00000000";
		ram_buffer(3495) := X"00000000";
		ram_buffer(3496) := X"00000000";
		ram_buffer(3497) := X"00000000";
		ram_buffer(3498) := X"00000000";
		ram_buffer(3499) := X"00000000";
		ram_buffer(3500) := X"00000000";
		ram_buffer(3501) := X"00000000";
		ram_buffer(3502) := X"00000000";
		ram_buffer(3503) := X"00000000";
		ram_buffer(3504) := X"00000000";
		ram_buffer(3505) := X"00000000";
		ram_buffer(3506) := X"00000000";
		ram_buffer(3507) := X"00000000";
		ram_buffer(3508) := X"00000000";
		ram_buffer(3509) := X"00000000";
		ram_buffer(3510) := X"00000000";
		ram_buffer(3511) := X"00000000";
		ram_buffer(3512) := X"00000000";
		ram_buffer(3513) := X"00000000";
		ram_buffer(3514) := X"00000000";
		ram_buffer(3515) := X"00000000";
		ram_buffer(3516) := X"00000000";
		ram_buffer(3517) := X"00000000";
		ram_buffer(3518) := X"00000000";
		ram_buffer(3519) := X"00000000";
		ram_buffer(3520) := X"00000000";
		ram_buffer(3521) := X"00000000";
		ram_buffer(3522) := X"00000000";
		ram_buffer(3523) := X"00000000";
		ram_buffer(3524) := X"00000000";
		ram_buffer(3525) := X"00000000";
		ram_buffer(3526) := X"00000000";
		ram_buffer(3527) := X"00000000";
		ram_buffer(3528) := X"00000000";
		ram_buffer(3529) := X"00000000";
		ram_buffer(3530) := X"00000000";
		ram_buffer(3531) := X"00000000";
		ram_buffer(3532) := X"00000000";
		ram_buffer(3533) := X"00000000";
		ram_buffer(3534) := X"00000000";
		ram_buffer(3535) := X"00000000";
		ram_buffer(3536) := X"00000000";
		ram_buffer(3537) := X"00000000";
		ram_buffer(3538) := X"00000000";
		ram_buffer(3539) := X"00000000";
		ram_buffer(3540) := X"00000000";
		ram_buffer(3541) := X"00000000";
		ram_buffer(3542) := X"00000000";
		ram_buffer(3543) := X"00000000";
		ram_buffer(3544) := X"00000000";
		ram_buffer(3545) := X"00000000";
		ram_buffer(3546) := X"00000000";
		ram_buffer(3547) := X"00000000";
		ram_buffer(3548) := X"00000000";
		ram_buffer(3549) := X"00000000";
		ram_buffer(3550) := X"00000000";
		ram_buffer(3551) := X"00000000";
		ram_buffer(3552) := X"00000000";
		ram_buffer(3553) := X"00000000";
		ram_buffer(3554) := X"00000000";
		ram_buffer(3555) := X"00000000";
		ram_buffer(3556) := X"00000000";
		ram_buffer(3557) := X"00000000";
		ram_buffer(3558) := X"00000000";
		ram_buffer(3559) := X"00000000";
		ram_buffer(3560) := X"00000000";
		ram_buffer(3561) := X"00000000";
		ram_buffer(3562) := X"00000000";
		ram_buffer(3563) := X"00000000";
		ram_buffer(3564) := X"00000000";
		ram_buffer(3565) := X"00000000";
		ram_buffer(3566) := X"00000000";
		ram_buffer(3567) := X"00000000";
		ram_buffer(3568) := X"00000000";
		ram_buffer(3569) := X"00000000";
		ram_buffer(3570) := X"00000000";
		ram_buffer(3571) := X"00000000";
		ram_buffer(3572) := X"00000000";
		ram_buffer(3573) := X"00000000";
		ram_buffer(3574) := X"00000000";
		ram_buffer(3575) := X"00000000";
		ram_buffer(3576) := X"00000000";
		ram_buffer(3577) := X"00000000";
		ram_buffer(3578) := X"00000000";
		ram_buffer(3579) := X"00000000";
		ram_buffer(3580) := X"00000000";
		ram_buffer(3581) := X"00000000";
		ram_buffer(3582) := X"00000000";
		ram_buffer(3583) := X"00000000";
		ram_buffer(3584) := X"00000000";
		ram_buffer(3585) := X"00000000";
		ram_buffer(3586) := X"00000000";
		ram_buffer(3587) := X"00000000";
		ram_buffer(3588) := X"00000000";
		ram_buffer(3589) := X"00000000";
		ram_buffer(3590) := X"00000000";
		ram_buffer(3591) := X"00000000";
		ram_buffer(3592) := X"00000000";
		ram_buffer(3593) := X"00000000";
		ram_buffer(3594) := X"00000000";
		ram_buffer(3595) := X"00000000";
		ram_buffer(3596) := X"00000000";
		ram_buffer(3597) := X"00000000";
		ram_buffer(3598) := X"00000000";
		ram_buffer(3599) := X"00000000";
		ram_buffer(3600) := X"00000000";
		ram_buffer(3601) := X"00000000";
		ram_buffer(3602) := X"00000000";
		ram_buffer(3603) := X"00000000";
		ram_buffer(3604) := X"00000000";
		ram_buffer(3605) := X"00000000";
		ram_buffer(3606) := X"00000000";
		ram_buffer(3607) := X"00000000";
		ram_buffer(3608) := X"00000000";
		ram_buffer(3609) := X"00000000";
		ram_buffer(3610) := X"00000000";
		ram_buffer(3611) := X"00000000";
		ram_buffer(3612) := X"00000000";
		ram_buffer(3613) := X"00000000";
		ram_buffer(3614) := X"00000000";
		ram_buffer(3615) := X"00000000";
		ram_buffer(3616) := X"00000000";
		ram_buffer(3617) := X"00000000";
		ram_buffer(3618) := X"00000000";
		ram_buffer(3619) := X"00000000";
		ram_buffer(3620) := X"00000000";
		ram_buffer(3621) := X"00000000";
		ram_buffer(3622) := X"00000000";
		ram_buffer(3623) := X"00000000";
		ram_buffer(3624) := X"00000000";
		ram_buffer(3625) := X"00000000";
		ram_buffer(3626) := X"00000000";
		ram_buffer(3627) := X"00000000";
		ram_buffer(3628) := X"00000000";
		ram_buffer(3629) := X"00000000";
		ram_buffer(3630) := X"00000000";
		ram_buffer(3631) := X"00000000";
		ram_buffer(3632) := X"00000000";
		ram_buffer(3633) := X"00000000";
		ram_buffer(3634) := X"00000000";
		ram_buffer(3635) := X"00000000";
		ram_buffer(3636) := X"00000000";
		ram_buffer(3637) := X"00000000";
		ram_buffer(3638) := X"00000000";
		ram_buffer(3639) := X"00000000";
		ram_buffer(3640) := X"00000000";
		ram_buffer(3641) := X"00000000";
		ram_buffer(3642) := X"00000000";
		ram_buffer(3643) := X"00000000";
		ram_buffer(3644) := X"00000000";
		ram_buffer(3645) := X"00000000";
		ram_buffer(3646) := X"00000000";
		ram_buffer(3647) := X"00000000";
		ram_buffer(3648) := X"00000000";
		ram_buffer(3649) := X"00000000";
		ram_buffer(3650) := X"00000000";
		ram_buffer(3651) := X"00000000";
		ram_buffer(3652) := X"00000000";
		ram_buffer(3653) := X"00000000";
		ram_buffer(3654) := X"00000000";
		ram_buffer(3655) := X"00000000";
		ram_buffer(3656) := X"00000000";
		ram_buffer(3657) := X"00000000";
		ram_buffer(3658) := X"00000000";
		ram_buffer(3659) := X"00000000";
		ram_buffer(3660) := X"00000000";
		ram_buffer(3661) := X"00000000";
		ram_buffer(3662) := X"00000000";
		ram_buffer(3663) := X"00000000";
		ram_buffer(3664) := X"00000000";
		ram_buffer(3665) := X"00000000";
		ram_buffer(3666) := X"00000000";
		ram_buffer(3667) := X"00000000";
		ram_buffer(3668) := X"00000000";
		ram_buffer(3669) := X"00000000";
		ram_buffer(3670) := X"00000000";
		ram_buffer(3671) := X"00000000";
		ram_buffer(3672) := X"00000000";
		ram_buffer(3673) := X"00000000";
		ram_buffer(3674) := X"00000000";
		ram_buffer(3675) := X"00000000";
		ram_buffer(3676) := X"00000000";
		ram_buffer(3677) := X"00000000";
		ram_buffer(3678) := X"00000000";
		ram_buffer(3679) := X"00000000";
		ram_buffer(3680) := X"00000000";
		ram_buffer(3681) := X"00000000";
		ram_buffer(3682) := X"00000000";
		ram_buffer(3683) := X"00000000";
		ram_buffer(3684) := X"00000000";
		ram_buffer(3685) := X"00000000";
		ram_buffer(3686) := X"00000000";
		ram_buffer(3687) := X"00000000";
		ram_buffer(3688) := X"00000000";
		ram_buffer(3689) := X"00000000";
		ram_buffer(3690) := X"00000000";
		ram_buffer(3691) := X"00000000";
		ram_buffer(3692) := X"00000000";
		ram_buffer(3693) := X"00000000";
		ram_buffer(3694) := X"00000000";
		ram_buffer(3695) := X"00000000";
		ram_buffer(3696) := X"00000000";
		ram_buffer(3697) := X"00000000";
		ram_buffer(3698) := X"00000000";
		ram_buffer(3699) := X"00000000";
		ram_buffer(3700) := X"00000000";
		ram_buffer(3701) := X"00000000";
		ram_buffer(3702) := X"00000000";
		ram_buffer(3703) := X"00000000";
		ram_buffer(3704) := X"00000000";
		ram_buffer(3705) := X"00000000";
		ram_buffer(3706) := X"00000000";
		ram_buffer(3707) := X"00000000";
		ram_buffer(3708) := X"00000000";
		ram_buffer(3709) := X"00000000";
		ram_buffer(3710) := X"00000000";
		ram_buffer(3711) := X"00000000";
		ram_buffer(3712) := X"00000000";
		ram_buffer(3713) := X"00000000";
		ram_buffer(3714) := X"00000000";
		ram_buffer(3715) := X"00000000";
		ram_buffer(3716) := X"00000000";
		ram_buffer(3717) := X"00000000";
		ram_buffer(3718) := X"00000000";
		ram_buffer(3719) := X"00000000";
		ram_buffer(3720) := X"00000000";
		ram_buffer(3721) := X"00000000";
		ram_buffer(3722) := X"00000000";
		ram_buffer(3723) := X"00000000";
		ram_buffer(3724) := X"00000000";
		ram_buffer(3725) := X"00000000";
		ram_buffer(3726) := X"00000000";
		ram_buffer(3727) := X"00000000";
		ram_buffer(3728) := X"00000000";
		ram_buffer(3729) := X"00000000";
		ram_buffer(3730) := X"00000000";
		ram_buffer(3731) := X"00000000";
		ram_buffer(3732) := X"00000000";
		ram_buffer(3733) := X"00000000";
		ram_buffer(3734) := X"00000000";
		ram_buffer(3735) := X"00000000";
		ram_buffer(3736) := X"00000000";
		ram_buffer(3737) := X"00000000";
		ram_buffer(3738) := X"00000000";
		ram_buffer(3739) := X"00000000";
		ram_buffer(3740) := X"00000000";
		ram_buffer(3741) := X"00000000";
		ram_buffer(3742) := X"00000000";
		ram_buffer(3743) := X"00000000";
		ram_buffer(3744) := X"00000000";
		ram_buffer(3745) := X"00000000";
		ram_buffer(3746) := X"00000000";
		ram_buffer(3747) := X"00000000";
		ram_buffer(3748) := X"00000000";
		ram_buffer(3749) := X"00000000";
		ram_buffer(3750) := X"00000000";
		ram_buffer(3751) := X"00000000";
		ram_buffer(3752) := X"00000000";
		ram_buffer(3753) := X"00000000";
		ram_buffer(3754) := X"00000000";
		ram_buffer(3755) := X"00000000";
		ram_buffer(3756) := X"00000000";
		ram_buffer(3757) := X"00000000";
		ram_buffer(3758) := X"00000000";
		ram_buffer(3759) := X"00000000";
		ram_buffer(3760) := X"00000000";
		ram_buffer(3761) := X"00000000";
		ram_buffer(3762) := X"00000000";
		ram_buffer(3763) := X"00000000";
		ram_buffer(3764) := X"00000000";
		ram_buffer(3765) := X"00000000";
		ram_buffer(3766) := X"00000000";
		ram_buffer(3767) := X"00000000";
		ram_buffer(3768) := X"00000000";
		ram_buffer(3769) := X"00000000";
		ram_buffer(3770) := X"00000000";
		ram_buffer(3771) := X"00000000";
		ram_buffer(3772) := X"00000000";
		ram_buffer(3773) := X"00000000";
		ram_buffer(3774) := X"00000000";
		ram_buffer(3775) := X"00000000";
		ram_buffer(3776) := X"00000000";
		ram_buffer(3777) := X"00000000";
		ram_buffer(3778) := X"00000000";
		ram_buffer(3779) := X"00000000";
		ram_buffer(3780) := X"00000000";
		ram_buffer(3781) := X"00000000";
		ram_buffer(3782) := X"00000000";
		ram_buffer(3783) := X"00000000";
		ram_buffer(3784) := X"00000000";
		ram_buffer(3785) := X"00000000";
		ram_buffer(3786) := X"00000000";
		ram_buffer(3787) := X"00000000";
		ram_buffer(3788) := X"00000000";
		ram_buffer(3789) := X"00000000";
		ram_buffer(3790) := X"00000000";
		ram_buffer(3791) := X"00000000";
		ram_buffer(3792) := X"00000000";
		ram_buffer(3793) := X"00000000";
		ram_buffer(3794) := X"00000000";
		ram_buffer(3795) := X"00000000";
		ram_buffer(3796) := X"00000000";
		ram_buffer(3797) := X"00000000";
		ram_buffer(3798) := X"00000000";
		ram_buffer(3799) := X"00000000";
		ram_buffer(3800) := X"00000000";
		ram_buffer(3801) := X"00000000";
		ram_buffer(3802) := X"00000000";
		ram_buffer(3803) := X"00000000";
		ram_buffer(3804) := X"00000000";
		ram_buffer(3805) := X"00000000";
		ram_buffer(3806) := X"00000000";
		ram_buffer(3807) := X"00000000";
		ram_buffer(3808) := X"00000000";
		ram_buffer(3809) := X"00000000";
		ram_buffer(3810) := X"00000000";
		ram_buffer(3811) := X"00000000";
		ram_buffer(3812) := X"00000000";
		ram_buffer(3813) := X"00000000";
		ram_buffer(3814) := X"00000000";
		ram_buffer(3815) := X"00000000";
		ram_buffer(3816) := X"00000000";
		ram_buffer(3817) := X"00000000";
		ram_buffer(3818) := X"00000000";
		ram_buffer(3819) := X"00000000";
		ram_buffer(3820) := X"00000000";
		ram_buffer(3821) := X"00000000";
		ram_buffer(3822) := X"00000000";
		ram_buffer(3823) := X"00000000";
		ram_buffer(3824) := X"00000000";
		ram_buffer(3825) := X"00000000";
		ram_buffer(3826) := X"00000000";
		ram_buffer(3827) := X"00000000";
		ram_buffer(3828) := X"00000000";
		ram_buffer(3829) := X"00000000";
		ram_buffer(3830) := X"00000000";
		ram_buffer(3831) := X"00000000";
		ram_buffer(3832) := X"00000000";
		ram_buffer(3833) := X"00000000";
		ram_buffer(3834) := X"00000000";
		ram_buffer(3835) := X"00000000";
		ram_buffer(3836) := X"00000000";
		ram_buffer(3837) := X"00000000";
		ram_buffer(3838) := X"00000000";
		ram_buffer(3839) := X"00000000";
		ram_buffer(3840) := X"00000000";
		ram_buffer(3841) := X"00000000";
		ram_buffer(3842) := X"00000000";
		ram_buffer(3843) := X"00000000";
		ram_buffer(3844) := X"00000000";
		ram_buffer(3845) := X"00000000";
		ram_buffer(3846) := X"00000000";
		ram_buffer(3847) := X"00000000";
		ram_buffer(3848) := X"00000000";
		ram_buffer(3849) := X"00000000";
		ram_buffer(3850) := X"00000000";
		ram_buffer(3851) := X"00000000";
		ram_buffer(3852) := X"00000000";
		ram_buffer(3853) := X"00000000";
		ram_buffer(3854) := X"00000000";
		ram_buffer(3855) := X"00000000";
		ram_buffer(3856) := X"00000000";
		ram_buffer(3857) := X"00000000";
		ram_buffer(3858) := X"00000000";
		ram_buffer(3859) := X"00000000";
		ram_buffer(3860) := X"00000000";
		ram_buffer(3861) := X"00000000";
		ram_buffer(3862) := X"00000000";
		ram_buffer(3863) := X"00000000";
		ram_buffer(3864) := X"00000000";
		ram_buffer(3865) := X"00000000";
		ram_buffer(3866) := X"00000000";
		ram_buffer(3867) := X"00000000";
		ram_buffer(3868) := X"00000000";
		ram_buffer(3869) := X"00000000";
		ram_buffer(3870) := X"00000000";
		ram_buffer(3871) := X"00000000";
		ram_buffer(3872) := X"00000000";
		ram_buffer(3873) := X"00000000";
		ram_buffer(3874) := X"00000000";
		ram_buffer(3875) := X"00000000";
		ram_buffer(3876) := X"00000000";
		ram_buffer(3877) := X"00000000";
		ram_buffer(3878) := X"00000000";
		ram_buffer(3879) := X"00000000";
		ram_buffer(3880) := X"00000000";
		ram_buffer(3881) := X"00000000";
		ram_buffer(3882) := X"00000000";
		ram_buffer(3883) := X"00000000";
		ram_buffer(3884) := X"00000000";
		ram_buffer(3885) := X"00000000";
		ram_buffer(3886) := X"00000000";
		ram_buffer(3887) := X"00000000";
		ram_buffer(3888) := X"00000000";
		ram_buffer(3889) := X"00000000";
		ram_buffer(3890) := X"00000000";
		ram_buffer(3891) := X"00000000";
		ram_buffer(3892) := X"00000000";
		ram_buffer(3893) := X"00000000";
		ram_buffer(3894) := X"00000000";
		ram_buffer(3895) := X"00000000";
		ram_buffer(3896) := X"00000000";
		ram_buffer(3897) := X"00000000";
		ram_buffer(3898) := X"00000000";
		ram_buffer(3899) := X"00000000";
		ram_buffer(3900) := X"00000000";
		ram_buffer(3901) := X"00000000";
		ram_buffer(3902) := X"00000000";
		ram_buffer(3903) := X"00000000";
		ram_buffer(3904) := X"00000000";
		ram_buffer(3905) := X"00000000";
		ram_buffer(3906) := X"00000000";
		ram_buffer(3907) := X"00000000";
		ram_buffer(3908) := X"00000000";
		ram_buffer(3909) := X"00000000";
		ram_buffer(3910) := X"00000000";
		ram_buffer(3911) := X"00000000";
		ram_buffer(3912) := X"00000000";
		ram_buffer(3913) := X"00000000";
		ram_buffer(3914) := X"00000000";
		ram_buffer(3915) := X"00000000";
		ram_buffer(3916) := X"00000000";
		ram_buffer(3917) := X"00000000";
		ram_buffer(3918) := X"00000000";
		ram_buffer(3919) := X"00000000";
		ram_buffer(3920) := X"00000000";
		ram_buffer(3921) := X"00000000";
		ram_buffer(3922) := X"00000000";
		ram_buffer(3923) := X"00000000";
		ram_buffer(3924) := X"00000000";
		ram_buffer(3925) := X"00000000";
		ram_buffer(3926) := X"00000000";
		ram_buffer(3927) := X"00000000";
		ram_buffer(3928) := X"00000000";
		ram_buffer(3929) := X"00000000";
		ram_buffer(3930) := X"00000000";
		ram_buffer(3931) := X"00000000";
		ram_buffer(3932) := X"00000000";
		ram_buffer(3933) := X"00000000";
		ram_buffer(3934) := X"00000000";
		ram_buffer(3935) := X"00000000";
		ram_buffer(3936) := X"00000000";
		ram_buffer(3937) := X"00000000";
		ram_buffer(3938) := X"00000000";
		ram_buffer(3939) := X"00000000";
		ram_buffer(3940) := X"00000000";
		ram_buffer(3941) := X"00000000";
		ram_buffer(3942) := X"00000000";
		ram_buffer(3943) := X"00000000";
		ram_buffer(3944) := X"00000000";
		ram_buffer(3945) := X"00000000";
		ram_buffer(3946) := X"00000000";
		ram_buffer(3947) := X"00000000";
		ram_buffer(3948) := X"00000000";
		ram_buffer(3949) := X"00000000";
		ram_buffer(3950) := X"00000000";
		ram_buffer(3951) := X"00000000";
		ram_buffer(3952) := X"00000000";
		ram_buffer(3953) := X"00000000";
		ram_buffer(3954) := X"00000000";
		ram_buffer(3955) := X"00000000";
		ram_buffer(3956) := X"00000000";
		ram_buffer(3957) := X"00000000";
		ram_buffer(3958) := X"00000000";
		ram_buffer(3959) := X"00000000";
		ram_buffer(3960) := X"00000000";
		ram_buffer(3961) := X"00000000";
		ram_buffer(3962) := X"00000000";
		ram_buffer(3963) := X"00000000";
		ram_buffer(3964) := X"00000000";
		ram_buffer(3965) := X"00000000";
		ram_buffer(3966) := X"00000000";
		ram_buffer(3967) := X"00000000";
		ram_buffer(3968) := X"00000000";
		ram_buffer(3969) := X"00000000";
		ram_buffer(3970) := X"00000000";
		ram_buffer(3971) := X"00000000";
		ram_buffer(3972) := X"00000000";
		ram_buffer(3973) := X"00000000";
		ram_buffer(3974) := X"00000000";
		ram_buffer(3975) := X"00000000";
		ram_buffer(3976) := X"00000000";
		ram_buffer(3977) := X"00000000";
		ram_buffer(3978) := X"00000000";
		ram_buffer(3979) := X"00000000";
		ram_buffer(3980) := X"00000000";
		ram_buffer(3981) := X"00000000";
		ram_buffer(3982) := X"00000000";
		ram_buffer(3983) := X"00000000";
		ram_buffer(3984) := X"00000000";
		ram_buffer(3985) := X"00000000";
		ram_buffer(3986) := X"00000000";
		ram_buffer(3987) := X"00000000";
		ram_buffer(3988) := X"00000000";
		ram_buffer(3989) := X"00000000";
		ram_buffer(3990) := X"00000000";
		ram_buffer(3991) := X"00000000";
		ram_buffer(3992) := X"00000000";
		ram_buffer(3993) := X"00000000";
		ram_buffer(3994) := X"00000000";
		ram_buffer(3995) := X"00000000";
		ram_buffer(3996) := X"00000000";
		ram_buffer(3997) := X"00000000";
		ram_buffer(3998) := X"00000000";
		ram_buffer(3999) := X"00000000";
		ram_buffer(4000) := X"00000000";
		ram_buffer(4001) := X"00000000";
		ram_buffer(4002) := X"00000000";
		ram_buffer(4003) := X"00000000";
		ram_buffer(4004) := X"00000000";
		ram_buffer(4005) := X"00000000";
		ram_buffer(4006) := X"00000000";
		ram_buffer(4007) := X"00000000";
		ram_buffer(4008) := X"00000000";
		ram_buffer(4009) := X"00000000";
		ram_buffer(4010) := X"00000000";
		ram_buffer(4011) := X"00000000";
		ram_buffer(4012) := X"00000000";
		ram_buffer(4013) := X"00000000";
		ram_buffer(4014) := X"00000000";
		ram_buffer(4015) := X"00000000";
		ram_buffer(4016) := X"00000000";
		ram_buffer(4017) := X"00000000";
		ram_buffer(4018) := X"00000000";
		ram_buffer(4019) := X"00000000";
		ram_buffer(4020) := X"00000000";
		ram_buffer(4021) := X"00000000";
		ram_buffer(4022) := X"00000000";
		ram_buffer(4023) := X"00000000";
		ram_buffer(4024) := X"00000000";
		ram_buffer(4025) := X"00000000";
		ram_buffer(4026) := X"00000000";
		ram_buffer(4027) := X"00000000";
		ram_buffer(4028) := X"00000000";
		ram_buffer(4029) := X"00000000";
		ram_buffer(4030) := X"00000000";
		ram_buffer(4031) := X"00000000";
		ram_buffer(4032) := X"00000000";
		ram_buffer(4033) := X"00000000";
		ram_buffer(4034) := X"00000000";
		ram_buffer(4035) := X"00000000";
		ram_buffer(4036) := X"00000000";
		ram_buffer(4037) := X"00000000";
		ram_buffer(4038) := X"00000000";
		ram_buffer(4039) := X"00000000";
		ram_buffer(4040) := X"00000000";
		ram_buffer(4041) := X"00000000";
		ram_buffer(4042) := X"00000000";
		ram_buffer(4043) := X"00000000";
		ram_buffer(4044) := X"00000000";
		ram_buffer(4045) := X"00000000";
		ram_buffer(4046) := X"00000000";
		ram_buffer(4047) := X"00000000";
		ram_buffer(4048) := X"00000000";
		ram_buffer(4049) := X"00000000";
		ram_buffer(4050) := X"00000000";
		ram_buffer(4051) := X"00000000";
		ram_buffer(4052) := X"00000000";
		ram_buffer(4053) := X"00000000";
		ram_buffer(4054) := X"00000000";
		ram_buffer(4055) := X"00000000";
		ram_buffer(4056) := X"00000000";
		ram_buffer(4057) := X"00000000";
		ram_buffer(4058) := X"00000000";
		ram_buffer(4059) := X"00000000";
		ram_buffer(4060) := X"00000000";
		ram_buffer(4061) := X"00000000";
		ram_buffer(4062) := X"00000000";
		ram_buffer(4063) := X"00000000";
		ram_buffer(4064) := X"00000000";
		ram_buffer(4065) := X"00000000";
		ram_buffer(4066) := X"00000000";
		ram_buffer(4067) := X"00000000";
		ram_buffer(4068) := X"00000000";
		ram_buffer(4069) := X"00000000";
		ram_buffer(4070) := X"00000000";
		ram_buffer(4071) := X"00000000";
		ram_buffer(4072) := X"00000000";
		ram_buffer(4073) := X"00000000";
		ram_buffer(4074) := X"00000000";
		ram_buffer(4075) := X"00000000";
		ram_buffer(4076) := X"00000000";
		ram_buffer(4077) := X"00000000";
		ram_buffer(4078) := X"00000000";
		ram_buffer(4079) := X"00000000";
		ram_buffer(4080) := X"00000000";
		ram_buffer(4081) := X"00000000";
		ram_buffer(4082) := X"00000000";
		ram_buffer(4083) := X"00000000";
		ram_buffer(4084) := X"00000000";
		ram_buffer(4085) := X"00000000";
		ram_buffer(4086) := X"00000000";
		ram_buffer(4087) := X"00000000";
		ram_buffer(4088) := X"00000000";
		ram_buffer(4089) := X"00000000";
		ram_buffer(4090) := X"00000000";
		ram_buffer(4091) := X"00000000";
		ram_buffer(4092) := X"00000000";
		ram_buffer(4093) := X"00000000";
		ram_buffer(4094) := X"00000000";
		ram_buffer(4095) := X"00000000";
		ram_buffer(4096) := X"00000000";
		ram_buffer(4097) := X"00000000";
		ram_buffer(4098) := X"00000000";
		ram_buffer(4099) := X"00000000";
		ram_buffer(4100) := X"00000000";
		ram_buffer(4101) := X"00000000";
		ram_buffer(4102) := X"00000000";
		ram_buffer(4103) := X"00000000";
		ram_buffer(4104) := X"00000000";
		ram_buffer(4105) := X"00000000";
		ram_buffer(4106) := X"00000000";
		ram_buffer(4107) := X"00000000";
		ram_buffer(4108) := X"00000000";
		ram_buffer(4109) := X"00000000";
		ram_buffer(4110) := X"00000000";
		ram_buffer(4111) := X"00000000";
		ram_buffer(4112) := X"00000000";
		ram_buffer(4113) := X"00000000";
		ram_buffer(4114) := X"00000000";
		ram_buffer(4115) := X"00000000";
		ram_buffer(4116) := X"00000000";
		ram_buffer(4117) := X"00000000";
		ram_buffer(4118) := X"00000000";
		ram_buffer(4119) := X"00000000";
		ram_buffer(4120) := X"00000000";
		ram_buffer(4121) := X"00000000";
		ram_buffer(4122) := X"00000000";
		ram_buffer(4123) := X"00000000";
		ram_buffer(4124) := X"00000000";
		ram_buffer(4125) := X"00000000";
		ram_buffer(4126) := X"00000000";
		ram_buffer(4127) := X"00000000";
		ram_buffer(4128) := X"00000000";
		ram_buffer(4129) := X"00000000";
		ram_buffer(4130) := X"00000000";
		ram_buffer(4131) := X"00000000";
		ram_buffer(4132) := X"00000000";
		ram_buffer(4133) := X"00000000";
		ram_buffer(4134) := X"00000000";
		ram_buffer(4135) := X"00000000";
		ram_buffer(4136) := X"00000000";
		ram_buffer(4137) := X"00000000";
		ram_buffer(4138) := X"00000000";
		ram_buffer(4139) := X"00000000";
		ram_buffer(4140) := X"00000000";
		ram_buffer(4141) := X"00000000";
		ram_buffer(4142) := X"00000000";
		ram_buffer(4143) := X"00000000";
		ram_buffer(4144) := X"00000000";
		ram_buffer(4145) := X"00000000";
		ram_buffer(4146) := X"00000000";
		ram_buffer(4147) := X"00000000";
		ram_buffer(4148) := X"00000000";
		ram_buffer(4149) := X"00000000";
		ram_buffer(4150) := X"00000000";
		ram_buffer(4151) := X"00000000";
		ram_buffer(4152) := X"00000000";
		ram_buffer(4153) := X"00000000";
		ram_buffer(4154) := X"00000000";
		ram_buffer(4155) := X"00000000";
		ram_buffer(4156) := X"00000000";
		ram_buffer(4157) := X"00000000";
		ram_buffer(4158) := X"00000000";
		ram_buffer(4159) := X"00000000";
		ram_buffer(4160) := X"00000000";
		ram_buffer(4161) := X"00000000";
		ram_buffer(4162) := X"00000000";
		ram_buffer(4163) := X"00000000";
		ram_buffer(4164) := X"00000000";
		ram_buffer(4165) := X"00000000";
		ram_buffer(4166) := X"00000000";
		ram_buffer(4167) := X"00000000";
		ram_buffer(4168) := X"00000000";
		ram_buffer(4169) := X"00000000";
		ram_buffer(4170) := X"00000000";
		ram_buffer(4171) := X"00000000";
		ram_buffer(4172) := X"00000000";
		ram_buffer(4173) := X"00000000";
		ram_buffer(4174) := X"00000000";
		ram_buffer(4175) := X"00000000";
		ram_buffer(4176) := X"00000000";
		ram_buffer(4177) := X"00000000";
		ram_buffer(4178) := X"00000000";
		ram_buffer(4179) := X"00000000";
		ram_buffer(4180) := X"00000000";
		ram_buffer(4181) := X"00000000";
		ram_buffer(4182) := X"00000000";
		ram_buffer(4183) := X"00000000";
		ram_buffer(4184) := X"00000000";
		ram_buffer(4185) := X"00000000";
		ram_buffer(4186) := X"00000000";
		ram_buffer(4187) := X"00000000";
		ram_buffer(4188) := X"00000000";
		ram_buffer(4189) := X"00000000";
		ram_buffer(4190) := X"00000000";
		ram_buffer(4191) := X"00000000";
		ram_buffer(4192) := X"00000000";
		ram_buffer(4193) := X"00000000";
		ram_buffer(4194) := X"00000000";
		ram_buffer(4195) := X"00000000";
		ram_buffer(4196) := X"00000000";
		ram_buffer(4197) := X"00000000";
		ram_buffer(4198) := X"00000000";
		ram_buffer(4199) := X"00000000";
		ram_buffer(4200) := X"00000000";
		ram_buffer(4201) := X"00000000";
		ram_buffer(4202) := X"00000000";
		ram_buffer(4203) := X"00000000";
		ram_buffer(4204) := X"00000000";
		ram_buffer(4205) := X"00000000";
		ram_buffer(4206) := X"00000000";
		ram_buffer(4207) := X"00000000";
		ram_buffer(4208) := X"00000000";
		ram_buffer(4209) := X"00000000";
		ram_buffer(4210) := X"00000000";
		ram_buffer(4211) := X"00000000";
		ram_buffer(4212) := X"00000000";
		ram_buffer(4213) := X"00000000";
		ram_buffer(4214) := X"00000000";
		ram_buffer(4215) := X"00000000";
		ram_buffer(4216) := X"00000000";
		ram_buffer(4217) := X"00000000";
		ram_buffer(4218) := X"00000000";
		ram_buffer(4219) := X"00000000";
		ram_buffer(4220) := X"00000000";
		ram_buffer(4221) := X"00000000";
		ram_buffer(4222) := X"00000000";
		ram_buffer(4223) := X"00000000";
		ram_buffer(4224) := X"00000000";
		ram_buffer(4225) := X"00000000";
		ram_buffer(4226) := X"00000000";
		ram_buffer(4227) := X"00000000";
		ram_buffer(4228) := X"00000000";
		ram_buffer(4229) := X"00000000";
		ram_buffer(4230) := X"00000000";
		ram_buffer(4231) := X"00000000";
		ram_buffer(4232) := X"00000000";
		ram_buffer(4233) := X"00000000";
		ram_buffer(4234) := X"00000000";
		ram_buffer(4235) := X"00000000";
		ram_buffer(4236) := X"00000000";
		ram_buffer(4237) := X"00000000";
		ram_buffer(4238) := X"00000000";
		ram_buffer(4239) := X"00000000";
		ram_buffer(4240) := X"00000000";
		ram_buffer(4241) := X"00000000";
		ram_buffer(4242) := X"00000000";
		ram_buffer(4243) := X"00000000";
		ram_buffer(4244) := X"00000000";
		ram_buffer(4245) := X"00000000";
		ram_buffer(4246) := X"00000000";
		ram_buffer(4247) := X"00000000";
		ram_buffer(4248) := X"00000000";
		ram_buffer(4249) := X"00000000";
		ram_buffer(4250) := X"00000000";
		ram_buffer(4251) := X"00000000";
		ram_buffer(4252) := X"00000000";
		ram_buffer(4253) := X"00000000";
		ram_buffer(4254) := X"00000000";
		ram_buffer(4255) := X"00000000";
		ram_buffer(4256) := X"00000000";
		ram_buffer(4257) := X"00000000";
		ram_buffer(4258) := X"00000000";
		ram_buffer(4259) := X"00000000";
		ram_buffer(4260) := X"00000000";
		ram_buffer(4261) := X"00000000";
		ram_buffer(4262) := X"00000000";
		ram_buffer(4263) := X"00000000";
		ram_buffer(4264) := X"00000000";
		ram_buffer(4265) := X"00000000";
		ram_buffer(4266) := X"00000000";
		ram_buffer(4267) := X"00000000";
		ram_buffer(4268) := X"00000000";
		ram_buffer(4269) := X"00000000";
		ram_buffer(4270) := X"00000000";
		ram_buffer(4271) := X"00000000";
		ram_buffer(4272) := X"00000000";
		ram_buffer(4273) := X"00000000";
		ram_buffer(4274) := X"00000000";
		ram_buffer(4275) := X"00000000";
		ram_buffer(4276) := X"00000000";
		ram_buffer(4277) := X"00000000";
		ram_buffer(4278) := X"00000000";
		ram_buffer(4279) := X"00000000";
		ram_buffer(4280) := X"00000000";
		ram_buffer(4281) := X"00000000";
		ram_buffer(4282) := X"00000000";
		ram_buffer(4283) := X"00000000";
		ram_buffer(4284) := X"00000000";
		ram_buffer(4285) := X"00000000";
		ram_buffer(4286) := X"00000000";
		ram_buffer(4287) := X"00000000";
		ram_buffer(4288) := X"00000000";
		ram_buffer(4289) := X"00000000";
		ram_buffer(4290) := X"00000000";
		ram_buffer(4291) := X"00000000";
		ram_buffer(4292) := X"00000000";
		ram_buffer(4293) := X"00000000";
		ram_buffer(4294) := X"00000000";
		ram_buffer(4295) := X"00000000";
		ram_buffer(4296) := X"00000000";
		ram_buffer(4297) := X"00000000";
		ram_buffer(4298) := X"00000000";
		ram_buffer(4299) := X"00000000";
		ram_buffer(4300) := X"00000000";
		ram_buffer(4301) := X"00000000";
		ram_buffer(4302) := X"00000000";
		ram_buffer(4303) := X"00000000";
		ram_buffer(4304) := X"00000000";
		ram_buffer(4305) := X"00000000";
		ram_buffer(4306) := X"00000000";
		ram_buffer(4307) := X"00000000";
		ram_buffer(4308) := X"00000000";
		ram_buffer(4309) := X"00000000";
		ram_buffer(4310) := X"00000000";
		ram_buffer(4311) := X"00000000";
		ram_buffer(4312) := X"00000000";
		ram_buffer(4313) := X"00000000";
		ram_buffer(4314) := X"00000000";
		ram_buffer(4315) := X"00000000";
		ram_buffer(4316) := X"00000000";
		ram_buffer(4317) := X"00000000";
		ram_buffer(4318) := X"00000000";
		ram_buffer(4319) := X"00000000";
		ram_buffer(4320) := X"00000000";
		ram_buffer(4321) := X"00000000";
		ram_buffer(4322) := X"00000000";
		ram_buffer(4323) := X"00000000";
		ram_buffer(4324) := X"00000000";
		ram_buffer(4325) := X"00000000";
		ram_buffer(4326) := X"00000000";
		ram_buffer(4327) := X"00000000";
		ram_buffer(4328) := X"00000000";
		ram_buffer(4329) := X"00000000";
		ram_buffer(4330) := X"00000000";
		ram_buffer(4331) := X"00000000";
		ram_buffer(4332) := X"00000000";
		ram_buffer(4333) := X"00000000";
		ram_buffer(4334) := X"00000000";
		ram_buffer(4335) := X"00000000";
		ram_buffer(4336) := X"00000000";
		ram_buffer(4337) := X"00000000";
		ram_buffer(4338) := X"00000000";
		ram_buffer(4339) := X"00000000";
		ram_buffer(4340) := X"00000000";
		ram_buffer(4341) := X"00000000";
		ram_buffer(4342) := X"00000000";
		ram_buffer(4343) := X"00000000";
		ram_buffer(4344) := X"00000000";
		ram_buffer(4345) := X"00000000";
		ram_buffer(4346) := X"00000000";
		ram_buffer(4347) := X"00000000";
		ram_buffer(4348) := X"00000000";
		ram_buffer(4349) := X"00000000";
		ram_buffer(4350) := X"00000000";
		ram_buffer(4351) := X"00000000";
		ram_buffer(4352) := X"00000000";
		ram_buffer(4353) := X"00000000";
		ram_buffer(4354) := X"00000000";
		ram_buffer(4355) := X"00000000";
		ram_buffer(4356) := X"00000000";
		ram_buffer(4357) := X"00000000";
		ram_buffer(4358) := X"00000000";
		ram_buffer(4359) := X"00000000";
		ram_buffer(4360) := X"00000000";
		ram_buffer(4361) := X"00000000";
		ram_buffer(4362) := X"00000000";
		ram_buffer(4363) := X"00000000";
		ram_buffer(4364) := X"00000000";
		ram_buffer(4365) := X"00000000";
		ram_buffer(4366) := X"00000000";
		ram_buffer(4367) := X"00000000";
		ram_buffer(4368) := X"00000000";
		ram_buffer(4369) := X"00000000";
		ram_buffer(4370) := X"00000000";
		ram_buffer(4371) := X"00000000";
		ram_buffer(4372) := X"00000000";
		ram_buffer(4373) := X"00000000";
		ram_buffer(4374) := X"00000000";
		ram_buffer(4375) := X"00000000";
		ram_buffer(4376) := X"00000000";
		ram_buffer(4377) := X"00000000";
		ram_buffer(4378) := X"00000000";
		ram_buffer(4379) := X"00000000";
		ram_buffer(4380) := X"00000000";
		ram_buffer(4381) := X"00000000";
		ram_buffer(4382) := X"00000000";
		ram_buffer(4383) := X"00000000";
		ram_buffer(4384) := X"00000000";
		ram_buffer(4385) := X"00000000";
		ram_buffer(4386) := X"00000000";
		ram_buffer(4387) := X"00000000";
		ram_buffer(4388) := X"00000000";
		ram_buffer(4389) := X"00000000";
		ram_buffer(4390) := X"00000000";
		ram_buffer(4391) := X"00000000";
		ram_buffer(4392) := X"00000000";
		ram_buffer(4393) := X"00000000";
		ram_buffer(4394) := X"00000000";
		ram_buffer(4395) := X"00000000";
		ram_buffer(4396) := X"00000000";
		ram_buffer(4397) := X"00000000";
		ram_buffer(4398) := X"00000000";
		ram_buffer(4399) := X"00000000";
		ram_buffer(4400) := X"00000000";
		ram_buffer(4401) := X"00000000";
		ram_buffer(4402) := X"00000000";
		ram_buffer(4403) := X"00000000";
		ram_buffer(4404) := X"00000000";
		ram_buffer(4405) := X"00000000";
		ram_buffer(4406) := X"00000000";
		ram_buffer(4407) := X"00000000";
		ram_buffer(4408) := X"00000000";
		ram_buffer(4409) := X"00000000";
		ram_buffer(4410) := X"00000000";
		ram_buffer(4411) := X"00000000";
		ram_buffer(4412) := X"00000000";
		ram_buffer(4413) := X"00000000";
		ram_buffer(4414) := X"00000000";
		ram_buffer(4415) := X"00000000";
		ram_buffer(4416) := X"00000000";
		ram_buffer(4417) := X"00000000";
		ram_buffer(4418) := X"00000000";
		ram_buffer(4419) := X"00000000";
		ram_buffer(4420) := X"00000000";
		ram_buffer(4421) := X"00000000";
		ram_buffer(4422) := X"00000000";
		ram_buffer(4423) := X"00000000";
		ram_buffer(4424) := X"00000000";
		ram_buffer(4425) := X"00000000";
		ram_buffer(4426) := X"00000000";
		ram_buffer(4427) := X"00000000";
		ram_buffer(4428) := X"00000000";
		ram_buffer(4429) := X"00000000";
		ram_buffer(4430) := X"00000000";
		ram_buffer(4431) := X"00000000";
		ram_buffer(4432) := X"00000000";
		ram_buffer(4433) := X"00000000";
		ram_buffer(4434) := X"00000000";
		ram_buffer(4435) := X"00000000";
		ram_buffer(4436) := X"00000000";
		ram_buffer(4437) := X"00000000";
		ram_buffer(4438) := X"00000000";
		ram_buffer(4439) := X"00000000";
		ram_buffer(4440) := X"00000000";
		ram_buffer(4441) := X"00000000";
		ram_buffer(4442) := X"00000000";
		ram_buffer(4443) := X"00000000";
		ram_buffer(4444) := X"00000000";
		ram_buffer(4445) := X"00000000";
		ram_buffer(4446) := X"00000000";
		ram_buffer(4447) := X"00000000";
		ram_buffer(4448) := X"00000000";
		ram_buffer(4449) := X"00000000";
		ram_buffer(4450) := X"00000000";
		ram_buffer(4451) := X"00000000";
		ram_buffer(4452) := X"00000000";
		ram_buffer(4453) := X"00000000";
		ram_buffer(4454) := X"00000000";
		ram_buffer(4455) := X"00000000";
		ram_buffer(4456) := X"00000000";
		ram_buffer(4457) := X"00000000";
		ram_buffer(4458) := X"00000000";
		ram_buffer(4459) := X"00000000";
		ram_buffer(4460) := X"00000000";
		ram_buffer(4461) := X"00000000";
		ram_buffer(4462) := X"00000000";
		ram_buffer(4463) := X"00000000";
		ram_buffer(4464) := X"00000000";
		ram_buffer(4465) := X"00000000";
		ram_buffer(4466) := X"00000000";
		ram_buffer(4467) := X"00000000";
		ram_buffer(4468) := X"00000000";
		ram_buffer(4469) := X"00000000";
		ram_buffer(4470) := X"00000000";
		ram_buffer(4471) := X"00000000";
		ram_buffer(4472) := X"00000000";
		ram_buffer(4473) := X"00000000";
		ram_buffer(4474) := X"00000000";
		ram_buffer(4475) := X"00000000";
		ram_buffer(4476) := X"00000000";
		ram_buffer(4477) := X"00000000";
		ram_buffer(4478) := X"00000000";
		ram_buffer(4479) := X"00000000";
		ram_buffer(4480) := X"00000000";
		ram_buffer(4481) := X"00000000";
		ram_buffer(4482) := X"00000000";
		ram_buffer(4483) := X"00000000";
		ram_buffer(4484) := X"00000000";
		ram_buffer(4485) := X"00000000";
		ram_buffer(4486) := X"00000000";
		ram_buffer(4487) := X"00000000";
		ram_buffer(4488) := X"00000000";
		ram_buffer(4489) := X"00000000";
		ram_buffer(4490) := X"00000000";
		ram_buffer(4491) := X"00000000";
		ram_buffer(4492) := X"00000000";
		ram_buffer(4493) := X"00000000";
		ram_buffer(4494) := X"00000000";
		ram_buffer(4495) := X"00000000";
		ram_buffer(4496) := X"00000000";
		ram_buffer(4497) := X"00000000";
		ram_buffer(4498) := X"00000000";
		ram_buffer(4499) := X"00000000";
		ram_buffer(4500) := X"00000000";
		ram_buffer(4501) := X"00000000";
		ram_buffer(4502) := X"00000000";
		ram_buffer(4503) := X"00000000";
		ram_buffer(4504) := X"00000000";
		ram_buffer(4505) := X"00000000";
		ram_buffer(4506) := X"00000000";
		ram_buffer(4507) := X"00000000";
		ram_buffer(4508) := X"00000000";
		ram_buffer(4509) := X"00000000";
		ram_buffer(4510) := X"00000000";
		ram_buffer(4511) := X"00000000";
		ram_buffer(4512) := X"00000000";
		ram_buffer(4513) := X"00000000";
		ram_buffer(4514) := X"00000000";
		ram_buffer(4515) := X"00000000";
		ram_buffer(4516) := X"00000000";
		ram_buffer(4517) := X"00000000";
		ram_buffer(4518) := X"00000000";
		ram_buffer(4519) := X"00000000";
		ram_buffer(4520) := X"00000000";
		ram_buffer(4521) := X"00000000";
		ram_buffer(4522) := X"00000000";
		ram_buffer(4523) := X"00000000";
		ram_buffer(4524) := X"00000000";
		ram_buffer(4525) := X"00000000";
		ram_buffer(4526) := X"00000000";
		ram_buffer(4527) := X"00000000";
		ram_buffer(4528) := X"00000000";
		ram_buffer(4529) := X"00000000";
		ram_buffer(4530) := X"00000000";
		ram_buffer(4531) := X"00000000";
		ram_buffer(4532) := X"00000000";
		ram_buffer(4533) := X"00000000";
		ram_buffer(4534) := X"00000000";
		ram_buffer(4535) := X"00000000";
		ram_buffer(4536) := X"00000000";
		ram_buffer(4537) := X"00000000";
		ram_buffer(4538) := X"00000000";
		ram_buffer(4539) := X"00000000";
		ram_buffer(4540) := X"00000000";
		ram_buffer(4541) := X"00000000";
		ram_buffer(4542) := X"00000000";
		ram_buffer(4543) := X"00000000";
		ram_buffer(4544) := X"00000000";
		ram_buffer(4545) := X"00000000";
		ram_buffer(4546) := X"00000000";
		ram_buffer(4547) := X"00000000";
		ram_buffer(4548) := X"00000000";
		ram_buffer(4549) := X"00000000";
		ram_buffer(4550) := X"00000000";
		ram_buffer(4551) := X"00000000";
		ram_buffer(4552) := X"00000000";
		ram_buffer(4553) := X"00000000";
		ram_buffer(4554) := X"00000000";
		ram_buffer(4555) := X"00000000";
		ram_buffer(4556) := X"00000000";
		ram_buffer(4557) := X"00000000";
		ram_buffer(4558) := X"00000000";
		ram_buffer(4559) := X"00000000";
		ram_buffer(4560) := X"00000000";
		ram_buffer(4561) := X"00000000";
		ram_buffer(4562) := X"00000000";
		ram_buffer(4563) := X"00000000";
		ram_buffer(4564) := X"00000000";
		ram_buffer(4565) := X"00000000";
		ram_buffer(4566) := X"00000000";
		ram_buffer(4567) := X"00000000";
		ram_buffer(4568) := X"00000000";
		ram_buffer(4569) := X"00000000";
		ram_buffer(4570) := X"00000000";
		ram_buffer(4571) := X"00000000";
		ram_buffer(4572) := X"00000000";
		ram_buffer(4573) := X"00000000";
		ram_buffer(4574) := X"00000000";
		ram_buffer(4575) := X"00000000";
		ram_buffer(4576) := X"00000000";
		ram_buffer(4577) := X"00000000";
		ram_buffer(4578) := X"00000000";
		ram_buffer(4579) := X"00000000";
		ram_buffer(4580) := X"00000000";
		ram_buffer(4581) := X"00000000";
		ram_buffer(4582) := X"00000000";
		ram_buffer(4583) := X"00000000";
		ram_buffer(4584) := X"00000000";
		ram_buffer(4585) := X"00000000";
		ram_buffer(4586) := X"00000000";
		ram_buffer(4587) := X"00000000";
		ram_buffer(4588) := X"00000000";
		ram_buffer(4589) := X"00000000";
		ram_buffer(4590) := X"00000000";
		ram_buffer(4591) := X"00000000";
		ram_buffer(4592) := X"00000000";
		ram_buffer(4593) := X"00000000";
		ram_buffer(4594) := X"00000000";
		ram_buffer(4595) := X"00000000";
		ram_buffer(4596) := X"00000000";
		ram_buffer(4597) := X"00000000";
		ram_buffer(4598) := X"00000000";
		ram_buffer(4599) := X"00000000";
		ram_buffer(4600) := X"00000000";
		ram_buffer(4601) := X"00000000";
		ram_buffer(4602) := X"00000000";
		ram_buffer(4603) := X"00000000";
		ram_buffer(4604) := X"00000000";
		ram_buffer(4605) := X"00000000";
		ram_buffer(4606) := X"00000000";
		ram_buffer(4607) := X"00000000";
		ram_buffer(4608) := X"00000000";
		ram_buffer(4609) := X"00000000";
		ram_buffer(4610) := X"00000000";
		ram_buffer(4611) := X"00000000";
		ram_buffer(4612) := X"00000000";
		ram_buffer(4613) := X"00000000";
		ram_buffer(4614) := X"00000000";
		ram_buffer(4615) := X"00000000";
		ram_buffer(4616) := X"00000000";
		ram_buffer(4617) := X"00000000";
		ram_buffer(4618) := X"00000000";
		ram_buffer(4619) := X"00000000";
		ram_buffer(4620) := X"00000000";
		ram_buffer(4621) := X"00000000";
		ram_buffer(4622) := X"00000000";
		ram_buffer(4623) := X"00000000";
		ram_buffer(4624) := X"00000000";
		ram_buffer(4625) := X"00000000";
		ram_buffer(4626) := X"00000000";
		ram_buffer(4627) := X"00000000";
		ram_buffer(4628) := X"00000000";
		ram_buffer(4629) := X"00000000";
		ram_buffer(4630) := X"00000000";
		ram_buffer(4631) := X"00000000";
		ram_buffer(4632) := X"00000000";
		ram_buffer(4633) := X"00000000";
		ram_buffer(4634) := X"00000000";
		ram_buffer(4635) := X"00000000";
		ram_buffer(4636) := X"00000000";
		ram_buffer(4637) := X"00000000";
		ram_buffer(4638) := X"00000000";
		ram_buffer(4639) := X"00000000";
		ram_buffer(4640) := X"00000000";
		ram_buffer(4641) := X"00000000";
		ram_buffer(4642) := X"00000000";
		ram_buffer(4643) := X"00000000";
		ram_buffer(4644) := X"00000000";
		ram_buffer(4645) := X"00000000";
		ram_buffer(4646) := X"00000000";
		ram_buffer(4647) := X"00000000";
		ram_buffer(4648) := X"00000000";
		ram_buffer(4649) := X"00000000";
		ram_buffer(4650) := X"00000000";
		ram_buffer(4651) := X"00000000";
		ram_buffer(4652) := X"00000000";
		ram_buffer(4653) := X"00000000";
		ram_buffer(4654) := X"00000000";
		ram_buffer(4655) := X"00000000";
		ram_buffer(4656) := X"00000000";
		ram_buffer(4657) := X"00000000";
		ram_buffer(4658) := X"00000000";
		ram_buffer(4659) := X"00000000";
		ram_buffer(4660) := X"00000000";
		ram_buffer(4661) := X"00000000";
		ram_buffer(4662) := X"00000000";
		ram_buffer(4663) := X"00000000";
		ram_buffer(4664) := X"00000000";
		ram_buffer(4665) := X"00000000";
		ram_buffer(4666) := X"00000000";
		ram_buffer(4667) := X"00000000";
		ram_buffer(4668) := X"00000000";
		ram_buffer(4669) := X"00000000";
		ram_buffer(4670) := X"00000000";
		ram_buffer(4671) := X"00000000";
		ram_buffer(4672) := X"00000000";
		ram_buffer(4673) := X"00000000";
		ram_buffer(4674) := X"00000000";
		ram_buffer(4675) := X"00000000";
		ram_buffer(4676) := X"00000000";
		ram_buffer(4677) := X"00000000";
		ram_buffer(4678) := X"00000000";
		ram_buffer(4679) := X"00000000";
		ram_buffer(4680) := X"00000000";
		ram_buffer(4681) := X"00000000";
		ram_buffer(4682) := X"00000000";
		ram_buffer(4683) := X"00000000";
		ram_buffer(4684) := X"00000000";
		ram_buffer(4685) := X"00000000";
		ram_buffer(4686) := X"00000000";
		ram_buffer(4687) := X"00000000";
		ram_buffer(4688) := X"00000000";
		ram_buffer(4689) := X"00000000";
		ram_buffer(4690) := X"00000000";
		ram_buffer(4691) := X"00000000";
		ram_buffer(4692) := X"00000000";
		ram_buffer(4693) := X"00000000";
		ram_buffer(4694) := X"00000000";
		ram_buffer(4695) := X"00000000";
		ram_buffer(4696) := X"00000000";
		ram_buffer(4697) := X"00000000";
		ram_buffer(4698) := X"00000000";
		ram_buffer(4699) := X"00000000";
		ram_buffer(4700) := X"00000000";
		ram_buffer(4701) := X"00000000";
		ram_buffer(4702) := X"00000000";
		ram_buffer(4703) := X"00000000";
		ram_buffer(4704) := X"00000000";
		ram_buffer(4705) := X"00000000";
		ram_buffer(4706) := X"00000000";
		ram_buffer(4707) := X"00000000";
		ram_buffer(4708) := X"00000000";
		ram_buffer(4709) := X"00000000";
		ram_buffer(4710) := X"00000000";
		ram_buffer(4711) := X"00000000";
		ram_buffer(4712) := X"00000000";
		ram_buffer(4713) := X"00000000";
		ram_buffer(4714) := X"00000000";
		ram_buffer(4715) := X"00000000";
		ram_buffer(4716) := X"00000000";
		ram_buffer(4717) := X"00000000";
		ram_buffer(4718) := X"00000000";
		ram_buffer(4719) := X"00000000";
		ram_buffer(4720) := X"00000000";
		ram_buffer(4721) := X"00000000";
		ram_buffer(4722) := X"00000000";
		ram_buffer(4723) := X"00000000";
		ram_buffer(4724) := X"00000000";
		ram_buffer(4725) := X"00000000";
		ram_buffer(4726) := X"00000000";
		ram_buffer(4727) := X"00000000";
		ram_buffer(4728) := X"00000000";
		ram_buffer(4729) := X"00000000";
		ram_buffer(4730) := X"00000000";
		ram_buffer(4731) := X"00000000";
		ram_buffer(4732) := X"00000000";
		ram_buffer(4733) := X"00000000";
		ram_buffer(4734) := X"00000000";
		ram_buffer(4735) := X"00000000";
		ram_buffer(4736) := X"00000000";
		ram_buffer(4737) := X"00000000";
		ram_buffer(4738) := X"00000000";
		ram_buffer(4739) := X"00000000";
		ram_buffer(4740) := X"00000000";
		ram_buffer(4741) := X"00000000";
		ram_buffer(4742) := X"00000000";
		ram_buffer(4743) := X"00000000";
		ram_buffer(4744) := X"00000000";
		ram_buffer(4745) := X"00000000";
		ram_buffer(4746) := X"00000000";
		ram_buffer(4747) := X"00000000";
		ram_buffer(4748) := X"00000000";
		ram_buffer(4749) := X"00000000";
		ram_buffer(4750) := X"00000000";
		ram_buffer(4751) := X"00000000";
		ram_buffer(4752) := X"00000000";
		ram_buffer(4753) := X"00000000";
		ram_buffer(4754) := X"00000000";
		ram_buffer(4755) := X"00000000";
		ram_buffer(4756) := X"00000000";
		ram_buffer(4757) := X"00000000";
		ram_buffer(4758) := X"00000000";
		ram_buffer(4759) := X"00000000";
		ram_buffer(4760) := X"00000000";
		ram_buffer(4761) := X"00000000";
		ram_buffer(4762) := X"00000000";
		ram_buffer(4763) := X"00000000";
		ram_buffer(4764) := X"00000000";
		ram_buffer(4765) := X"00000000";
		ram_buffer(4766) := X"00000000";
		ram_buffer(4767) := X"00000000";
		ram_buffer(4768) := X"00000000";
		ram_buffer(4769) := X"00000000";
		ram_buffer(4770) := X"00000000";
		ram_buffer(4771) := X"00000000";
		ram_buffer(4772) := X"00000000";
		ram_buffer(4773) := X"00000000";
		ram_buffer(4774) := X"00000000";
		ram_buffer(4775) := X"00000000";
		ram_buffer(4776) := X"00000000";
		ram_buffer(4777) := X"00000000";
		ram_buffer(4778) := X"00000000";
		ram_buffer(4779) := X"00000000";
		ram_buffer(4780) := X"00000000";
		ram_buffer(4781) := X"00000000";
		ram_buffer(4782) := X"00000000";
		ram_buffer(4783) := X"00000000";
		ram_buffer(4784) := X"00000000";
		ram_buffer(4785) := X"00000000";
		ram_buffer(4786) := X"00000000";
		ram_buffer(4787) := X"00000000";
		ram_buffer(4788) := X"00000000";
		ram_buffer(4789) := X"00000000";
		ram_buffer(4790) := X"00000000";
		ram_buffer(4791) := X"00000000";
		ram_buffer(4792) := X"00000000";
		ram_buffer(4793) := X"00000000";
		ram_buffer(4794) := X"00000000";
		ram_buffer(4795) := X"00000000";
		ram_buffer(4796) := X"00000000";
		ram_buffer(4797) := X"00000000";
		ram_buffer(4798) := X"00000000";
		ram_buffer(4799) := X"00000000";
		ram_buffer(4800) := X"00000000";
		ram_buffer(4801) := X"00000000";
		ram_buffer(4802) := X"00000000";
		ram_buffer(4803) := X"00000000";
		ram_buffer(4804) := X"00000000";
		ram_buffer(4805) := X"00000000";
		ram_buffer(4806) := X"00000000";
		ram_buffer(4807) := X"00000000";
		ram_buffer(4808) := X"00000000";
		ram_buffer(4809) := X"00000000";
		ram_buffer(4810) := X"00000000";
		ram_buffer(4811) := X"00000000";
		ram_buffer(4812) := X"00000000";
		ram_buffer(4813) := X"00000000";
		ram_buffer(4814) := X"00000000";
		ram_buffer(4815) := X"00000000";
		ram_buffer(4816) := X"00000000";
		ram_buffer(4817) := X"00000000";
		ram_buffer(4818) := X"00000000";
		ram_buffer(4819) := X"00000000";
		ram_buffer(4820) := X"00000000";
		ram_buffer(4821) := X"00000000";
		ram_buffer(4822) := X"00000000";
		ram_buffer(4823) := X"00000000";
		ram_buffer(4824) := X"00000000";
		ram_buffer(4825) := X"00000000";
		ram_buffer(4826) := X"00000000";
		ram_buffer(4827) := X"00000000";
		ram_buffer(4828) := X"00000000";
		ram_buffer(4829) := X"00000000";
		ram_buffer(4830) := X"00000000";
		ram_buffer(4831) := X"00000000";
		ram_buffer(4832) := X"00000000";
		ram_buffer(4833) := X"00000000";
		ram_buffer(4834) := X"00000000";
		ram_buffer(4835) := X"00000000";
		ram_buffer(4836) := X"00000000";
		ram_buffer(4837) := X"00000000";
		ram_buffer(4838) := X"00000000";
		ram_buffer(4839) := X"00000000";
		ram_buffer(4840) := X"00000000";
		ram_buffer(4841) := X"00000000";
		ram_buffer(4842) := X"00000000";
		ram_buffer(4843) := X"00000000";
		ram_buffer(4844) := X"00000000";
		ram_buffer(4845) := X"00000000";
		ram_buffer(4846) := X"00000000";
		ram_buffer(4847) := X"00000000";
		ram_buffer(4848) := X"00000000";
		ram_buffer(4849) := X"00000000";
		ram_buffer(4850) := X"00000000";
		ram_buffer(4851) := X"00000000";
		ram_buffer(4852) := X"00000000";
		ram_buffer(4853) := X"00000000";
		ram_buffer(4854) := X"00000000";
		ram_buffer(4855) := X"00000000";
		ram_buffer(4856) := X"00000000";
		ram_buffer(4857) := X"00000000";
		ram_buffer(4858) := X"00000000";
		ram_buffer(4859) := X"00000000";
		ram_buffer(4860) := X"00000000";
		ram_buffer(4861) := X"00000000";
		ram_buffer(4862) := X"00000000";
		ram_buffer(4863) := X"00000000";
		ram_buffer(4864) := X"00000000";
		ram_buffer(4865) := X"00000000";
		ram_buffer(4866) := X"00000000";
		ram_buffer(4867) := X"00000000";
		ram_buffer(4868) := X"00000000";
		ram_buffer(4869) := X"00000000";
		ram_buffer(4870) := X"00000000";
		ram_buffer(4871) := X"00000000";
		ram_buffer(4872) := X"00000000";
		ram_buffer(4873) := X"00000000";
		ram_buffer(4874) := X"00000000";
		ram_buffer(4875) := X"00000000";
		ram_buffer(4876) := X"00000000";
		ram_buffer(4877) := X"00000000";
		ram_buffer(4878) := X"00000000";
		ram_buffer(4879) := X"00000000";
		ram_buffer(4880) := X"00000000";
		ram_buffer(4881) := X"00000000";
		ram_buffer(4882) := X"00000000";
		ram_buffer(4883) := X"00000000";
		ram_buffer(4884) := X"00000000";
		ram_buffer(4885) := X"00000000";
		ram_buffer(4886) := X"00000000";
		ram_buffer(4887) := X"00000000";
		ram_buffer(4888) := X"00000000";
		ram_buffer(4889) := X"00000000";
		ram_buffer(4890) := X"00000000";
		ram_buffer(4891) := X"00000000";
		ram_buffer(4892) := X"00000000";
		ram_buffer(4893) := X"00000000";
		ram_buffer(4894) := X"00000000";
		ram_buffer(4895) := X"00000000";
		ram_buffer(4896) := X"00000000";
		ram_buffer(4897) := X"00000000";
		ram_buffer(4898) := X"00000000";
		ram_buffer(4899) := X"00000000";
		ram_buffer(4900) := X"00000000";
		ram_buffer(4901) := X"00000000";
		ram_buffer(4902) := X"00000000";
		ram_buffer(4903) := X"00000000";
		ram_buffer(4904) := X"00000000";
		ram_buffer(4905) := X"00000000";
		ram_buffer(4906) := X"00000000";
		ram_buffer(4907) := X"00000000";
		ram_buffer(4908) := X"00000000";
		ram_buffer(4909) := X"00000000";
		ram_buffer(4910) := X"00000000";
		ram_buffer(4911) := X"00000000";
		ram_buffer(4912) := X"00000000";
		ram_buffer(4913) := X"00000000";
		ram_buffer(4914) := X"00000000";
		ram_buffer(4915) := X"00000000";
		ram_buffer(4916) := X"00000000";
		ram_buffer(4917) := X"00000000";
		ram_buffer(4918) := X"00000000";
		ram_buffer(4919) := X"00000000";
		ram_buffer(4920) := X"00000000";
		ram_buffer(4921) := X"00000000";
		ram_buffer(4922) := X"00000000";
		ram_buffer(4923) := X"00000000";
		ram_buffer(4924) := X"00000000";
		ram_buffer(4925) := X"00000000";
		ram_buffer(4926) := X"00000000";
		ram_buffer(4927) := X"00000000";
		ram_buffer(4928) := X"00000000";
		ram_buffer(4929) := X"00000000";
		ram_buffer(4930) := X"00000000";
		ram_buffer(4931) := X"00000000";
		ram_buffer(4932) := X"00000000";
		ram_buffer(4933) := X"00000000";
		ram_buffer(4934) := X"00000000";
		ram_buffer(4935) := X"00000000";
		ram_buffer(4936) := X"00000000";
		ram_buffer(4937) := X"00000000";
		ram_buffer(4938) := X"00000000";
		ram_buffer(4939) := X"00000000";
		ram_buffer(4940) := X"00000000";
		ram_buffer(4941) := X"00000000";
		ram_buffer(4942) := X"00000000";
		ram_buffer(4943) := X"00000000";
		ram_buffer(4944) := X"00000000";
		ram_buffer(4945) := X"00000000";
		ram_buffer(4946) := X"00000000";
		ram_buffer(4947) := X"00000000";
		ram_buffer(4948) := X"00000000";
		ram_buffer(4949) := X"00000000";
		ram_buffer(4950) := X"00000000";
		ram_buffer(4951) := X"00000000";
		ram_buffer(4952) := X"00000000";
		ram_buffer(4953) := X"00000000";
		ram_buffer(4954) := X"00000000";
		ram_buffer(4955) := X"00000000";
		ram_buffer(4956) := X"00000000";
		ram_buffer(4957) := X"00000000";
		ram_buffer(4958) := X"00000000";
		ram_buffer(4959) := X"00000000";
		ram_buffer(4960) := X"00000000";
		ram_buffer(4961) := X"00000000";
		ram_buffer(4962) := X"00000000";
		ram_buffer(4963) := X"00000000";
		ram_buffer(4964) := X"00000000";
		ram_buffer(4965) := X"00000000";
		ram_buffer(4966) := X"00000000";
		ram_buffer(4967) := X"00000000";
		ram_buffer(4968) := X"00000000";
		ram_buffer(4969) := X"00000000";
		ram_buffer(4970) := X"00000000";
		ram_buffer(4971) := X"00000000";
		ram_buffer(4972) := X"00000000";
		ram_buffer(4973) := X"00000000";
		ram_buffer(4974) := X"00000000";
		ram_buffer(4975) := X"00000000";
		ram_buffer(4976) := X"00000000";
		ram_buffer(4977) := X"00000000";
		ram_buffer(4978) := X"00000000";
		ram_buffer(4979) := X"00000000";
		ram_buffer(4980) := X"00000000";
		ram_buffer(4981) := X"00000000";
		ram_buffer(4982) := X"00000000";
		ram_buffer(4983) := X"00000000";
		ram_buffer(4984) := X"00000000";
		ram_buffer(4985) := X"00000000";
		ram_buffer(4986) := X"00000000";
		ram_buffer(4987) := X"00000000";
		ram_buffer(4988) := X"00000000";
		ram_buffer(4989) := X"00000000";
		ram_buffer(4990) := X"00000000";
		ram_buffer(4991) := X"00000000";
		ram_buffer(4992) := X"00000000";
		ram_buffer(4993) := X"00000000";
		ram_buffer(4994) := X"00000000";
		ram_buffer(4995) := X"00000000";
		ram_buffer(4996) := X"00000000";
		ram_buffer(4997) := X"00000000";
		ram_buffer(4998) := X"00000000";
		ram_buffer(4999) := X"00000000";
		ram_buffer(5000) := X"00000000";
		ram_buffer(5001) := X"00000000";
		ram_buffer(5002) := X"00000000";
		ram_buffer(5003) := X"00000000";
		ram_buffer(5004) := X"00000000";
		ram_buffer(5005) := X"00000000";
		ram_buffer(5006) := X"00000000";
		ram_buffer(5007) := X"00000000";
		ram_buffer(5008) := X"00000000";
		ram_buffer(5009) := X"00000000";
		ram_buffer(5010) := X"00000000";
		ram_buffer(5011) := X"00000000";
		ram_buffer(5012) := X"00000000";
		ram_buffer(5013) := X"00000000";
		ram_buffer(5014) := X"00000000";
		ram_buffer(5015) := X"00000000";
		ram_buffer(5016) := X"00000000";
		ram_buffer(5017) := X"00000000";
		ram_buffer(5018) := X"00000000";
		ram_buffer(5019) := X"00000000";
		ram_buffer(5020) := X"00000000";
		ram_buffer(5021) := X"00000000";
		ram_buffer(5022) := X"00000000";
		ram_buffer(5023) := X"00000000";
		ram_buffer(5024) := X"00000000";
		ram_buffer(5025) := X"00000000";
		ram_buffer(5026) := X"00000000";
		ram_buffer(5027) := X"00000000";
		ram_buffer(5028) := X"00000000";
		ram_buffer(5029) := X"00000000";
		ram_buffer(5030) := X"00000000";
		ram_buffer(5031) := X"00000000";
		ram_buffer(5032) := X"00000000";
		ram_buffer(5033) := X"00000000";
		ram_buffer(5034) := X"00000000";
		ram_buffer(5035) := X"00000000";
		ram_buffer(5036) := X"00000000";
		ram_buffer(5037) := X"00000000";
		ram_buffer(5038) := X"00000000";
		ram_buffer(5039) := X"00000000";
		ram_buffer(5040) := X"00000000";
		ram_buffer(5041) := X"00000000";
		ram_buffer(5042) := X"00000000";
		ram_buffer(5043) := X"00000000";
		ram_buffer(5044) := X"00000000";
		ram_buffer(5045) := X"00000000";
		ram_buffer(5046) := X"00000000";
		ram_buffer(5047) := X"00000000";
		ram_buffer(5048) := X"00000000";
		ram_buffer(5049) := X"00000000";
		ram_buffer(5050) := X"00000000";
		ram_buffer(5051) := X"00000000";
		ram_buffer(5052) := X"00000000";
		ram_buffer(5053) := X"00000000";
		ram_buffer(5054) := X"00000000";
		ram_buffer(5055) := X"00000000";
		ram_buffer(5056) := X"00000000";
		ram_buffer(5057) := X"00000000";
		ram_buffer(5058) := X"00000000";
		ram_buffer(5059) := X"00000000";
		ram_buffer(5060) := X"00000000";
		ram_buffer(5061) := X"00000000";
		ram_buffer(5062) := X"00000000";
		ram_buffer(5063) := X"00000000";
		ram_buffer(5064) := X"00000000";
		ram_buffer(5065) := X"00000000";
		ram_buffer(5066) := X"00000000";
		ram_buffer(5067) := X"00000000";
		ram_buffer(5068) := X"00000000";
		ram_buffer(5069) := X"00000000";
		ram_buffer(5070) := X"00000000";
		ram_buffer(5071) := X"00000000";
		ram_buffer(5072) := X"00000000";
		ram_buffer(5073) := X"00000000";
		ram_buffer(5074) := X"00000000";
		ram_buffer(5075) := X"00000000";
		ram_buffer(5076) := X"00000000";
		ram_buffer(5077) := X"00000000";
		ram_buffer(5078) := X"00000000";
		ram_buffer(5079) := X"00000000";
		ram_buffer(5080) := X"00000000";
		ram_buffer(5081) := X"00000000";
		ram_buffer(5082) := X"00000000";
		ram_buffer(5083) := X"00000000";
		ram_buffer(5084) := X"00000000";
		ram_buffer(5085) := X"00000000";
		ram_buffer(5086) := X"00000000";
		ram_buffer(5087) := X"00000000";
		ram_buffer(5088) := X"00000000";
		ram_buffer(5089) := X"00000000";
		ram_buffer(5090) := X"00000000";
		ram_buffer(5091) := X"00000000";
		ram_buffer(5092) := X"00000000";
		ram_buffer(5093) := X"00000000";
		ram_buffer(5094) := X"00000000";
		ram_buffer(5095) := X"00000000";
		ram_buffer(5096) := X"00000000";
		ram_buffer(5097) := X"00000000";
		ram_buffer(5098) := X"00000000";
		ram_buffer(5099) := X"00000000";
		ram_buffer(5100) := X"00000000";
		ram_buffer(5101) := X"00000000";
		ram_buffer(5102) := X"00000000";
		ram_buffer(5103) := X"00000000";
		ram_buffer(5104) := X"00000000";
		ram_buffer(5105) := X"00000000";
		ram_buffer(5106) := X"00000000";
		ram_buffer(5107) := X"00000000";
		ram_buffer(5108) := X"00000000";
		ram_buffer(5109) := X"00000000";
		ram_buffer(5110) := X"00000000";
		ram_buffer(5111) := X"00000000";
		ram_buffer(5112) := X"00000000";
		ram_buffer(5113) := X"00000000";
		ram_buffer(5114) := X"00000000";
		ram_buffer(5115) := X"00000000";
		ram_buffer(5116) := X"00000000";
		ram_buffer(5117) := X"00000000";
		ram_buffer(5118) := X"00000000";
		ram_buffer(5119) := X"00000000";
		ram_buffer(5120) := X"00000000";
		ram_buffer(5121) := X"00000000";
		ram_buffer(5122) := X"00000000";
		ram_buffer(5123) := X"00000000";
		ram_buffer(5124) := X"00000000";
		ram_buffer(5125) := X"00000000";
		ram_buffer(5126) := X"00000000";
		ram_buffer(5127) := X"00000000";
		ram_buffer(5128) := X"00000000";
		ram_buffer(5129) := X"00000000";
		ram_buffer(5130) := X"00000000";
		ram_buffer(5131) := X"00000000";
		ram_buffer(5132) := X"00000000";
		ram_buffer(5133) := X"00000000";
		ram_buffer(5134) := X"00000000";
		ram_buffer(5135) := X"00000000";
		ram_buffer(5136) := X"00000000";
		ram_buffer(5137) := X"00000000";
		ram_buffer(5138) := X"00000000";
		ram_buffer(5139) := X"00000000";
		ram_buffer(5140) := X"00000000";
		ram_buffer(5141) := X"00000000";
		ram_buffer(5142) := X"00000000";
		ram_buffer(5143) := X"00000000";
		ram_buffer(5144) := X"00000000";
		ram_buffer(5145) := X"00000000";
		ram_buffer(5146) := X"00000000";
		ram_buffer(5147) := X"00000000";
		ram_buffer(5148) := X"00000000";
		ram_buffer(5149) := X"00000000";
		ram_buffer(5150) := X"00000000";
		ram_buffer(5151) := X"00000000";
		ram_buffer(5152) := X"00000000";
		ram_buffer(5153) := X"00000000";
		ram_buffer(5154) := X"00000000";
		ram_buffer(5155) := X"00000000";
		ram_buffer(5156) := X"00000000";
		ram_buffer(5157) := X"00000000";
		ram_buffer(5158) := X"00000000";
		ram_buffer(5159) := X"00000000";
		ram_buffer(5160) := X"00000000";
		ram_buffer(5161) := X"00000000";
		ram_buffer(5162) := X"00000000";
		ram_buffer(5163) := X"00000000";
		ram_buffer(5164) := X"00000000";
		ram_buffer(5165) := X"00000000";
		ram_buffer(5166) := X"00000000";
		ram_buffer(5167) := X"00000000";
		ram_buffer(5168) := X"00000000";
		ram_buffer(5169) := X"00000000";
		ram_buffer(5170) := X"00000000";
		ram_buffer(5171) := X"00000000";
		ram_buffer(5172) := X"00000000";
		ram_buffer(5173) := X"00000000";
		ram_buffer(5174) := X"00000000";
		ram_buffer(5175) := X"00000000";
		ram_buffer(5176) := X"00000000";
		ram_buffer(5177) := X"00000000";
		ram_buffer(5178) := X"00000000";
		ram_buffer(5179) := X"00000000";
		ram_buffer(5180) := X"00000000";
		ram_buffer(5181) := X"00000000";
		ram_buffer(5182) := X"00000000";
		ram_buffer(5183) := X"00000000";
		ram_buffer(5184) := X"00000000";
		ram_buffer(5185) := X"00000000";
		ram_buffer(5186) := X"00000000";
		ram_buffer(5187) := X"00000000";
		ram_buffer(5188) := X"00000000";
		ram_buffer(5189) := X"00000000";
		ram_buffer(5190) := X"00000000";
		ram_buffer(5191) := X"00000000";
		ram_buffer(5192) := X"00000000";
		ram_buffer(5193) := X"00000000";
		ram_buffer(5194) := X"00000000";
		ram_buffer(5195) := X"00000000";
		ram_buffer(5196) := X"00000000";
		ram_buffer(5197) := X"00000000";
		ram_buffer(5198) := X"00000000";
		ram_buffer(5199) := X"00000000";
		ram_buffer(5200) := X"00000000";
		ram_buffer(5201) := X"00000000";
		ram_buffer(5202) := X"00000000";
		ram_buffer(5203) := X"00000000";
		ram_buffer(5204) := X"00000000";
		ram_buffer(5205) := X"00000000";
		ram_buffer(5206) := X"00000000";
		ram_buffer(5207) := X"00000000";
		ram_buffer(5208) := X"00000000";
		ram_buffer(5209) := X"00000000";
		ram_buffer(5210) := X"00000000";
		ram_buffer(5211) := X"00000000";
		ram_buffer(5212) := X"00000000";
		ram_buffer(5213) := X"00000000";
		ram_buffer(5214) := X"00000000";
		ram_buffer(5215) := X"00000000";
		ram_buffer(5216) := X"00000000";
		ram_buffer(5217) := X"00000000";
		ram_buffer(5218) := X"00000000";
		ram_buffer(5219) := X"00000000";
		ram_buffer(5220) := X"00000000";
		ram_buffer(5221) := X"00000000";
		ram_buffer(5222) := X"00000000";
		ram_buffer(5223) := X"00000000";
		ram_buffer(5224) := X"00000000";
		ram_buffer(5225) := X"00000000";
		ram_buffer(5226) := X"00000000";
		ram_buffer(5227) := X"00000000";
		ram_buffer(5228) := X"00000000";
		ram_buffer(5229) := X"00000000";
		ram_buffer(5230) := X"00000000";
		ram_buffer(5231) := X"00000000";
		ram_buffer(5232) := X"00000000";
		ram_buffer(5233) := X"00000000";
		ram_buffer(5234) := X"00000000";
		ram_buffer(5235) := X"00000000";
		ram_buffer(5236) := X"00000000";
		ram_buffer(5237) := X"00000000";
		ram_buffer(5238) := X"00000000";
		ram_buffer(5239) := X"00000000";
		ram_buffer(5240) := X"00000000";
		ram_buffer(5241) := X"00000000";
		ram_buffer(5242) := X"00000000";
		ram_buffer(5243) := X"00000000";
		ram_buffer(5244) := X"00000000";
		ram_buffer(5245) := X"00000000";
		ram_buffer(5246) := X"00000000";
		ram_buffer(5247) := X"00000000";
		ram_buffer(5248) := X"00000000";
		ram_buffer(5249) := X"00000000";
		ram_buffer(5250) := X"00000000";
		ram_buffer(5251) := X"00000000";
		ram_buffer(5252) := X"00000000";
		ram_buffer(5253) := X"00000000";
		ram_buffer(5254) := X"00000000";
		ram_buffer(5255) := X"00000000";
		ram_buffer(5256) := X"00000000";
		ram_buffer(5257) := X"00000000";
		ram_buffer(5258) := X"00000000";
		ram_buffer(5259) := X"00000000";
		ram_buffer(5260) := X"00000000";
		ram_buffer(5261) := X"00000000";
		ram_buffer(5262) := X"00000000";
		ram_buffer(5263) := X"00000000";
		ram_buffer(5264) := X"00000000";
		ram_buffer(5265) := X"00000000";
		ram_buffer(5266) := X"00000000";
		ram_buffer(5267) := X"00000000";
		ram_buffer(5268) := X"00000000";
		ram_buffer(5269) := X"00000000";
		ram_buffer(5270) := X"00000000";
		ram_buffer(5271) := X"00000000";
		ram_buffer(5272) := X"00000000";
		ram_buffer(5273) := X"00000000";
		ram_buffer(5274) := X"00000000";
		ram_buffer(5275) := X"00000000";
		ram_buffer(5276) := X"00000000";
		ram_buffer(5277) := X"00000000";
		ram_buffer(5278) := X"00000000";
		ram_buffer(5279) := X"00000000";
		ram_buffer(5280) := X"00000000";
		ram_buffer(5281) := X"00000000";
		ram_buffer(5282) := X"00000000";
		ram_buffer(5283) := X"00000000";
		ram_buffer(5284) := X"00000000";
		ram_buffer(5285) := X"00000000";
		ram_buffer(5286) := X"00000000";
		ram_buffer(5287) := X"00000000";
		ram_buffer(5288) := X"00000000";
		ram_buffer(5289) := X"00000000";
		ram_buffer(5290) := X"00000000";
		ram_buffer(5291) := X"00000000";
		ram_buffer(5292) := X"00000000";
		ram_buffer(5293) := X"00000000";
		ram_buffer(5294) := X"00000000";
		ram_buffer(5295) := X"00000000";
		ram_buffer(5296) := X"00000000";
		ram_buffer(5297) := X"00000000";
		ram_buffer(5298) := X"00000000";
		ram_buffer(5299) := X"00000000";
		ram_buffer(5300) := X"00000000";
		ram_buffer(5301) := X"00000000";
		ram_buffer(5302) := X"00000000";
		ram_buffer(5303) := X"00000000";
		ram_buffer(5304) := X"00000000";
		ram_buffer(5305) := X"00000000";
		ram_buffer(5306) := X"00000000";
		ram_buffer(5307) := X"00000000";
		ram_buffer(5308) := X"00000000";
		ram_buffer(5309) := X"00000000";
		ram_buffer(5310) := X"00000000";
		ram_buffer(5311) := X"00000000";
		ram_buffer(5312) := X"00000000";
		ram_buffer(5313) := X"00000000";
		ram_buffer(5314) := X"00000000";
		ram_buffer(5315) := X"00000000";
		ram_buffer(5316) := X"00000000";
		ram_buffer(5317) := X"00000000";
		ram_buffer(5318) := X"00000000";
		ram_buffer(5319) := X"00000000";
		ram_buffer(5320) := X"00000000";
		ram_buffer(5321) := X"00000000";
		ram_buffer(5322) := X"00000000";
		ram_buffer(5323) := X"00000000";
		ram_buffer(5324) := X"00000000";
		ram_buffer(5325) := X"00000000";
		ram_buffer(5326) := X"00000000";
		ram_buffer(5327) := X"00000000";
		ram_buffer(5328) := X"00000000";
		ram_buffer(5329) := X"00000000";
		ram_buffer(5330) := X"00000000";
		ram_buffer(5331) := X"00000000";
		ram_buffer(5332) := X"00000000";
		ram_buffer(5333) := X"00000000";
		ram_buffer(5334) := X"00000000";
		ram_buffer(5335) := X"00000000";
		ram_buffer(5336) := X"00000000";
		ram_buffer(5337) := X"00000000";
		ram_buffer(5338) := X"00000000";
		ram_buffer(5339) := X"00000000";
		ram_buffer(5340) := X"00000000";
		ram_buffer(5341) := X"00000000";
		ram_buffer(5342) := X"00000000";
		ram_buffer(5343) := X"00000000";
		ram_buffer(5344) := X"00000000";
		ram_buffer(5345) := X"00000000";
		ram_buffer(5346) := X"00000000";
		ram_buffer(5347) := X"00000000";
		ram_buffer(5348) := X"00000000";
		ram_buffer(5349) := X"00000000";
		ram_buffer(5350) := X"00000000";
		ram_buffer(5351) := X"00000000";
		ram_buffer(5352) := X"00000000";
		ram_buffer(5353) := X"00000000";
		ram_buffer(5354) := X"00000000";
		ram_buffer(5355) := X"00000000";
		ram_buffer(5356) := X"00000000";
		ram_buffer(5357) := X"00000000";
		ram_buffer(5358) := X"00000000";
		ram_buffer(5359) := X"00000000";
		ram_buffer(5360) := X"00000000";
		ram_buffer(5361) := X"00000000";
		ram_buffer(5362) := X"00000000";
		ram_buffer(5363) := X"00000000";
		ram_buffer(5364) := X"00000000";
		ram_buffer(5365) := X"00000000";
		ram_buffer(5366) := X"00000000";
		ram_buffer(5367) := X"00000000";
		ram_buffer(5368) := X"00000000";
		ram_buffer(5369) := X"00000000";
		ram_buffer(5370) := X"00000000";
		ram_buffer(5371) := X"00000000";
		ram_buffer(5372) := X"00000000";
		ram_buffer(5373) := X"00000000";
		ram_buffer(5374) := X"00000000";
		ram_buffer(5375) := X"00000000";
		ram_buffer(5376) := X"00000000";
		ram_buffer(5377) := X"00000000";
		ram_buffer(5378) := X"00000000";
		ram_buffer(5379) := X"00000000";
		ram_buffer(5380) := X"00000000";
		ram_buffer(5381) := X"00000000";
		ram_buffer(5382) := X"00000000";
		ram_buffer(5383) := X"00000000";
		ram_buffer(5384) := X"00000000";
		ram_buffer(5385) := X"00000000";
		ram_buffer(5386) := X"00000000";
		ram_buffer(5387) := X"00000000";
		ram_buffer(5388) := X"00000000";
		ram_buffer(5389) := X"00000000";
		ram_buffer(5390) := X"00000000";
		ram_buffer(5391) := X"00000000";
		ram_buffer(5392) := X"00000000";
		ram_buffer(5393) := X"00000000";
		ram_buffer(5394) := X"00000000";
		ram_buffer(5395) := X"00000000";
		ram_buffer(5396) := X"00000000";
		ram_buffer(5397) := X"00000000";
		ram_buffer(5398) := X"00000000";
		ram_buffer(5399) := X"00000000";
		ram_buffer(5400) := X"00000000";
		ram_buffer(5401) := X"00000000";
		ram_buffer(5402) := X"00000000";
		ram_buffer(5403) := X"00000000";
		ram_buffer(5404) := X"00000000";
		ram_buffer(5405) := X"00000000";
		ram_buffer(5406) := X"00000000";
		ram_buffer(5407) := X"00000000";
		ram_buffer(5408) := X"00000000";
		ram_buffer(5409) := X"00000000";
		ram_buffer(5410) := X"00000000";
		ram_buffer(5411) := X"00000000";
		ram_buffer(5412) := X"00000000";
		ram_buffer(5413) := X"00000000";
		ram_buffer(5414) := X"00000000";
		ram_buffer(5415) := X"00000000";
		ram_buffer(5416) := X"00000000";
		ram_buffer(5417) := X"00000000";
		ram_buffer(5418) := X"00000000";
		ram_buffer(5419) := X"00000000";
		ram_buffer(5420) := X"00000000";
		ram_buffer(5421) := X"00000000";
		ram_buffer(5422) := X"00000000";
		ram_buffer(5423) := X"00000000";
		ram_buffer(5424) := X"00000000";
		ram_buffer(5425) := X"00000000";
		ram_buffer(5426) := X"00000000";
		ram_buffer(5427) := X"00000000";
		ram_buffer(5428) := X"00000000";
		ram_buffer(5429) := X"00000000";
		ram_buffer(5430) := X"00000000";
		ram_buffer(5431) := X"00000000";
		ram_buffer(5432) := X"00000000";
		ram_buffer(5433) := X"00000000";
		ram_buffer(5434) := X"00000000";
		ram_buffer(5435) := X"00000000";
		ram_buffer(5436) := X"00000000";
		ram_buffer(5437) := X"00000000";
		ram_buffer(5438) := X"00000000";
		ram_buffer(5439) := X"00000000";
		ram_buffer(5440) := X"00000000";
		ram_buffer(5441) := X"00000000";
		ram_buffer(5442) := X"00000000";
		ram_buffer(5443) := X"00000000";
		ram_buffer(5444) := X"00000000";
		ram_buffer(5445) := X"00000000";
		ram_buffer(5446) := X"00000000";
		ram_buffer(5447) := X"00000000";
		ram_buffer(5448) := X"00000000";
		ram_buffer(5449) := X"00000000";
		ram_buffer(5450) := X"00000000";
		ram_buffer(5451) := X"00000000";
		ram_buffer(5452) := X"00000000";
		ram_buffer(5453) := X"00000000";
		ram_buffer(5454) := X"00000000";
		ram_buffer(5455) := X"00000000";
		ram_buffer(5456) := X"00000000";
		ram_buffer(5457) := X"00000000";
		ram_buffer(5458) := X"00000000";
		ram_buffer(5459) := X"00000000";
		ram_buffer(5460) := X"00000000";
		ram_buffer(5461) := X"00000000";
		ram_buffer(5462) := X"00000000";
		ram_buffer(5463) := X"00000000";
		ram_buffer(5464) := X"00000000";
		ram_buffer(5465) := X"00000000";
		ram_buffer(5466) := X"00000000";
		ram_buffer(5467) := X"00000000";
		ram_buffer(5468) := X"00000000";
		ram_buffer(5469) := X"00000000";
		ram_buffer(5470) := X"00000000";
		ram_buffer(5471) := X"00000000";
		ram_buffer(5472) := X"00000000";
		ram_buffer(5473) := X"00000000";
		ram_buffer(5474) := X"00000000";
		ram_buffer(5475) := X"00000000";
		ram_buffer(5476) := X"00000000";
		ram_buffer(5477) := X"00000000";
		ram_buffer(5478) := X"00000000";
		ram_buffer(5479) := X"00000000";
		ram_buffer(5480) := X"00000000";
		ram_buffer(5481) := X"00000000";
		ram_buffer(5482) := X"00000000";
		ram_buffer(5483) := X"00000000";
		ram_buffer(5484) := X"00000000";
		ram_buffer(5485) := X"00000000";
		ram_buffer(5486) := X"00000000";
		ram_buffer(5487) := X"00000000";
		ram_buffer(5488) := X"00000000";
		ram_buffer(5489) := X"00000000";
		ram_buffer(5490) := X"00000000";
		ram_buffer(5491) := X"00000000";
		ram_buffer(5492) := X"00000000";
		ram_buffer(5493) := X"00000000";
		ram_buffer(5494) := X"00000000";
		ram_buffer(5495) := X"00000000";
		ram_buffer(5496) := X"00000000";
		ram_buffer(5497) := X"00000000";
		ram_buffer(5498) := X"00000000";
		ram_buffer(5499) := X"00000000";
		ram_buffer(5500) := X"00000000";
		ram_buffer(5501) := X"00000000";
		ram_buffer(5502) := X"00000000";
		ram_buffer(5503) := X"00000000";
		ram_buffer(5504) := X"00000000";
		ram_buffer(5505) := X"00000000";
		ram_buffer(5506) := X"00000000";
		ram_buffer(5507) := X"00000000";
		ram_buffer(5508) := X"00000000";
		ram_buffer(5509) := X"00000000";
		ram_buffer(5510) := X"00000000";
		ram_buffer(5511) := X"00000000";
		ram_buffer(5512) := X"00000000";
		ram_buffer(5513) := X"00000000";
		ram_buffer(5514) := X"00000000";
		ram_buffer(5515) := X"00000000";
		ram_buffer(5516) := X"00000000";
		ram_buffer(5517) := X"00000000";
		ram_buffer(5518) := X"00000000";
		ram_buffer(5519) := X"00000000";
		ram_buffer(5520) := X"00000000";
		ram_buffer(5521) := X"00000000";
		ram_buffer(5522) := X"00000000";
		ram_buffer(5523) := X"00000000";
		ram_buffer(5524) := X"00000000";
		ram_buffer(5525) := X"00000000";
		ram_buffer(5526) := X"00000000";
		ram_buffer(5527) := X"00000000";
		ram_buffer(5528) := X"00000000";
		ram_buffer(5529) := X"00000000";
		ram_buffer(5530) := X"00000000";
		ram_buffer(5531) := X"00000000";
		ram_buffer(5532) := X"00000000";
		ram_buffer(5533) := X"00000000";
		ram_buffer(5534) := X"00000000";
		ram_buffer(5535) := X"00000000";
		ram_buffer(5536) := X"00000000";
		ram_buffer(5537) := X"00000000";
		ram_buffer(5538) := X"00000000";
		ram_buffer(5539) := X"00000000";
		ram_buffer(5540) := X"00000000";
		ram_buffer(5541) := X"00000000";
		ram_buffer(5542) := X"00000000";
		ram_buffer(5543) := X"00000000";
		ram_buffer(5544) := X"00000000";
		ram_buffer(5545) := X"00000000";
		ram_buffer(5546) := X"00000000";
		ram_buffer(5547) := X"00000000";
		ram_buffer(5548) := X"00000000";
		ram_buffer(5549) := X"00000000";
		ram_buffer(5550) := X"00000000";
		ram_buffer(5551) := X"00000000";
		ram_buffer(5552) := X"00000000";
		ram_buffer(5553) := X"00000000";
		ram_buffer(5554) := X"00000000";
		ram_buffer(5555) := X"00000000";
		ram_buffer(5556) := X"00000000";
		ram_buffer(5557) := X"00000000";
		ram_buffer(5558) := X"00000000";
		ram_buffer(5559) := X"00000000";
		ram_buffer(5560) := X"00000000";
		ram_buffer(5561) := X"00000000";
		ram_buffer(5562) := X"00000000";
		ram_buffer(5563) := X"00000000";
		ram_buffer(5564) := X"00000000";
		ram_buffer(5565) := X"00000000";
		ram_buffer(5566) := X"00000000";
		ram_buffer(5567) := X"00000000";
		ram_buffer(5568) := X"00000000";
		ram_buffer(5569) := X"00000000";
		ram_buffer(5570) := X"00000000";
		ram_buffer(5571) := X"00000000";
		ram_buffer(5572) := X"00000000";
		ram_buffer(5573) := X"00000000";
		ram_buffer(5574) := X"00000000";
		ram_buffer(5575) := X"00000000";
		ram_buffer(5576) := X"00000000";
		ram_buffer(5577) := X"00000000";
		ram_buffer(5578) := X"00000000";
		ram_buffer(5579) := X"00000000";
		ram_buffer(5580) := X"00000000";
		ram_buffer(5581) := X"00000000";
		ram_buffer(5582) := X"00000000";
		ram_buffer(5583) := X"00000000";
		ram_buffer(5584) := X"00000000";
		ram_buffer(5585) := X"00000000";
		ram_buffer(5586) := X"00000000";
		ram_buffer(5587) := X"00000000";
		ram_buffer(5588) := X"00000000";
		ram_buffer(5589) := X"00000000";
		ram_buffer(5590) := X"00000000";
		ram_buffer(5591) := X"00000000";
		ram_buffer(5592) := X"00000000";
		ram_buffer(5593) := X"00000000";
		ram_buffer(5594) := X"00000000";
		ram_buffer(5595) := X"00000000";
		ram_buffer(5596) := X"00000000";
		ram_buffer(5597) := X"00000000";
		ram_buffer(5598) := X"00000000";
		ram_buffer(5599) := X"00000000";
		ram_buffer(5600) := X"00000000";
		ram_buffer(5601) := X"00000000";
		ram_buffer(5602) := X"00000000";
		ram_buffer(5603) := X"00000000";
		ram_buffer(5604) := X"00000000";
		ram_buffer(5605) := X"00000000";
		ram_buffer(5606) := X"00000000";
		ram_buffer(5607) := X"00000000";
		ram_buffer(5608) := X"00000000";
		ram_buffer(5609) := X"00000000";
		ram_buffer(5610) := X"00000000";
		ram_buffer(5611) := X"00000000";
		ram_buffer(5612) := X"00000000";
		ram_buffer(5613) := X"00000000";
		ram_buffer(5614) := X"00000000";
		ram_buffer(5615) := X"00000000";
		ram_buffer(5616) := X"00000000";
		ram_buffer(5617) := X"00000000";
		ram_buffer(5618) := X"00000000";
		ram_buffer(5619) := X"00000000";
		ram_buffer(5620) := X"00000000";
		ram_buffer(5621) := X"00000000";
		ram_buffer(5622) := X"00000000";
		ram_buffer(5623) := X"00000000";
		ram_buffer(5624) := X"00000000";
		ram_buffer(5625) := X"00000000";
		ram_buffer(5626) := X"00000000";
		ram_buffer(5627) := X"00000000";
		ram_buffer(5628) := X"00000000";
		ram_buffer(5629) := X"00000000";
		ram_buffer(5630) := X"00000000";
		ram_buffer(5631) := X"00000000";
		ram_buffer(5632) := X"00000000";
		ram_buffer(5633) := X"00000000";
		ram_buffer(5634) := X"00000000";
		ram_buffer(5635) := X"00000000";
		ram_buffer(5636) := X"00000000";
		ram_buffer(5637) := X"00000000";
		ram_buffer(5638) := X"00000000";
		ram_buffer(5639) := X"00000000";
		ram_buffer(5640) := X"00000000";
		ram_buffer(5641) := X"00000000";
		ram_buffer(5642) := X"00000000";
		ram_buffer(5643) := X"00000000";
		ram_buffer(5644) := X"00000000";
		ram_buffer(5645) := X"00000000";
		ram_buffer(5646) := X"00000000";
		ram_buffer(5647) := X"00000000";
		ram_buffer(5648) := X"00000000";
		ram_buffer(5649) := X"00000000";
		ram_buffer(5650) := X"00000000";
		ram_buffer(5651) := X"00000000";
		ram_buffer(5652) := X"00000000";
		ram_buffer(5653) := X"00000000";
		ram_buffer(5654) := X"00000000";
		ram_buffer(5655) := X"00000000";
		ram_buffer(5656) := X"00000000";
		ram_buffer(5657) := X"00000000";
		ram_buffer(5658) := X"00000000";
		ram_buffer(5659) := X"00000000";
		ram_buffer(5660) := X"00000000";
		ram_buffer(5661) := X"00000000";
		ram_buffer(5662) := X"00000000";
		ram_buffer(5663) := X"00000000";
		ram_buffer(5664) := X"00000000";
		ram_buffer(5665) := X"00000000";
		ram_buffer(5666) := X"00000000";
		ram_buffer(5667) := X"00000000";
		ram_buffer(5668) := X"00000000";
		ram_buffer(5669) := X"00000000";
		ram_buffer(5670) := X"00000000";
		ram_buffer(5671) := X"00000000";
		ram_buffer(5672) := X"00000000";
		ram_buffer(5673) := X"00000000";
		ram_buffer(5674) := X"00000000";
		ram_buffer(5675) := X"00000000";
		ram_buffer(5676) := X"00000000";
		ram_buffer(5677) := X"00000000";
		ram_buffer(5678) := X"00000000";
		ram_buffer(5679) := X"00000000";
		ram_buffer(5680) := X"00000000";
		ram_buffer(5681) := X"00000000";
		ram_buffer(5682) := X"00000000";
		ram_buffer(5683) := X"00000000";
		ram_buffer(5684) := X"00000000";
		ram_buffer(5685) := X"00000000";
		ram_buffer(5686) := X"00000000";
		ram_buffer(5687) := X"00000000";
		ram_buffer(5688) := X"00000000";
		ram_buffer(5689) := X"00000000";
		ram_buffer(5690) := X"00000000";
		ram_buffer(5691) := X"00000000";
		ram_buffer(5692) := X"00000000";
		ram_buffer(5693) := X"00000000";
		ram_buffer(5694) := X"00000000";
		ram_buffer(5695) := X"00000000";
		ram_buffer(5696) := X"00000000";
		ram_buffer(5697) := X"00000000";
		ram_buffer(5698) := X"00000000";
		ram_buffer(5699) := X"00000000";
		ram_buffer(5700) := X"00000000";
		ram_buffer(5701) := X"00000000";
		ram_buffer(5702) := X"00000000";
		ram_buffer(5703) := X"00000000";
		ram_buffer(5704) := X"00000000";
		ram_buffer(5705) := X"00000000";
		ram_buffer(5706) := X"00000000";
		ram_buffer(5707) := X"00000000";
		ram_buffer(5708) := X"00000000";
		ram_buffer(5709) := X"00000000";
		ram_buffer(5710) := X"00000000";
		ram_buffer(5711) := X"00000000";
		ram_buffer(5712) := X"00000000";
		ram_buffer(5713) := X"00000000";
		ram_buffer(5714) := X"00000000";
		ram_buffer(5715) := X"00000000";
		ram_buffer(5716) := X"00000000";
		ram_buffer(5717) := X"00000000";
		ram_buffer(5718) := X"00000000";
		ram_buffer(5719) := X"00000000";
		ram_buffer(5720) := X"00000000";
		ram_buffer(5721) := X"00000000";
		ram_buffer(5722) := X"00000000";
		ram_buffer(5723) := X"00000000";
		ram_buffer(5724) := X"00000000";
		ram_buffer(5725) := X"00000000";
		ram_buffer(5726) := X"00000000";
		ram_buffer(5727) := X"00000000";
		ram_buffer(5728) := X"00000000";
		ram_buffer(5729) := X"00000000";
		ram_buffer(5730) := X"00000000";
		ram_buffer(5731) := X"00000000";
		ram_buffer(5732) := X"00000000";
		ram_buffer(5733) := X"00000000";
		ram_buffer(5734) := X"00000000";
		ram_buffer(5735) := X"00000000";
		ram_buffer(5736) := X"00000000";
		ram_buffer(5737) := X"00000000";
		ram_buffer(5738) := X"00000000";
		ram_buffer(5739) := X"00000000";
		ram_buffer(5740) := X"00000000";
		ram_buffer(5741) := X"00000000";
		ram_buffer(5742) := X"00000000";
		ram_buffer(5743) := X"00000000";
		ram_buffer(5744) := X"00000000";
		ram_buffer(5745) := X"00000000";
		ram_buffer(5746) := X"00000000";
		ram_buffer(5747) := X"00000000";
		ram_buffer(5748) := X"00000000";
		ram_buffer(5749) := X"00000000";
		ram_buffer(5750) := X"00000000";
		ram_buffer(5751) := X"00000000";
		ram_buffer(5752) := X"00000000";
		ram_buffer(5753) := X"00000000";
		ram_buffer(5754) := X"00000000";
		ram_buffer(5755) := X"00000000";
		ram_buffer(5756) := X"00000000";
		ram_buffer(5757) := X"00000000";
		ram_buffer(5758) := X"00000000";
		ram_buffer(5759) := X"00000000";
		ram_buffer(5760) := X"00000000";
		ram_buffer(5761) := X"00000000";
		ram_buffer(5762) := X"00000000";
		ram_buffer(5763) := X"00000000";
		ram_buffer(5764) := X"00000000";
		ram_buffer(5765) := X"00000000";
		ram_buffer(5766) := X"00000000";
		ram_buffer(5767) := X"00000000";
		ram_buffer(5768) := X"00000000";
		ram_buffer(5769) := X"00000000";
		ram_buffer(5770) := X"00000000";
		ram_buffer(5771) := X"00000000";
		ram_buffer(5772) := X"00000000";
		ram_buffer(5773) := X"00000000";
		ram_buffer(5774) := X"00000000";
		ram_buffer(5775) := X"00000000";
		ram_buffer(5776) := X"00000000";
		ram_buffer(5777) := X"00000000";
		ram_buffer(5778) := X"00000000";
		ram_buffer(5779) := X"00000000";
		ram_buffer(5780) := X"00000000";
		ram_buffer(5781) := X"00000000";
		ram_buffer(5782) := X"00000000";
		ram_buffer(5783) := X"00000000";
		ram_buffer(5784) := X"00000000";
		ram_buffer(5785) := X"00000000";
		ram_buffer(5786) := X"00000000";
		ram_buffer(5787) := X"00000000";
		ram_buffer(5788) := X"00000000";
		ram_buffer(5789) := X"00000000";
		ram_buffer(5790) := X"00000000";
		ram_buffer(5791) := X"00000000";
		ram_buffer(5792) := X"00000000";
		ram_buffer(5793) := X"00000000";
		ram_buffer(5794) := X"00000000";
		ram_buffer(5795) := X"00000000";
		ram_buffer(5796) := X"00000000";
		ram_buffer(5797) := X"00000000";
		ram_buffer(5798) := X"00000000";
		ram_buffer(5799) := X"00000000";
		ram_buffer(5800) := X"00000000";
		ram_buffer(5801) := X"00000000";
		ram_buffer(5802) := X"00000000";
		ram_buffer(5803) := X"00000000";
		ram_buffer(5804) := X"00000000";
		ram_buffer(5805) := X"00000000";
		ram_buffer(5806) := X"00000000";
		ram_buffer(5807) := X"00000000";
		ram_buffer(5808) := X"00000000";
		ram_buffer(5809) := X"00000000";
		ram_buffer(5810) := X"00000000";
		ram_buffer(5811) := X"00000000";
		ram_buffer(5812) := X"00000000";
		ram_buffer(5813) := X"00000000";
		ram_buffer(5814) := X"00000000";
		ram_buffer(5815) := X"00000000";
		ram_buffer(5816) := X"00000000";
		ram_buffer(5817) := X"00000000";
		ram_buffer(5818) := X"00000000";
		ram_buffer(5819) := X"00000000";
		ram_buffer(5820) := X"00000000";
		ram_buffer(5821) := X"00000000";
		ram_buffer(5822) := X"00000000";
		ram_buffer(5823) := X"00000000";
		ram_buffer(5824) := X"00000000";
		ram_buffer(5825) := X"00000000";
		ram_buffer(5826) := X"00000000";
		ram_buffer(5827) := X"00000000";
		ram_buffer(5828) := X"00000000";
		ram_buffer(5829) := X"00000000";
		ram_buffer(5830) := X"00000000";
		ram_buffer(5831) := X"00000000";
		ram_buffer(5832) := X"00000000";
		ram_buffer(5833) := X"00000000";
		ram_buffer(5834) := X"00000000";
		ram_buffer(5835) := X"00000000";
		ram_buffer(5836) := X"00000000";
		ram_buffer(5837) := X"00000000";
		ram_buffer(5838) := X"00000000";
		ram_buffer(5839) := X"00000000";
		ram_buffer(5840) := X"00000000";
		ram_buffer(5841) := X"00000000";
		ram_buffer(5842) := X"00000000";
		ram_buffer(5843) := X"00000000";
		ram_buffer(5844) := X"00000000";
		ram_buffer(5845) := X"00000000";
		ram_buffer(5846) := X"00000000";
		ram_buffer(5847) := X"00000000";
		ram_buffer(5848) := X"00000000";
		ram_buffer(5849) := X"00000000";
		ram_buffer(5850) := X"00000000";
		ram_buffer(5851) := X"00000000";
		ram_buffer(5852) := X"00000000";
		ram_buffer(5853) := X"00000000";
		ram_buffer(5854) := X"00000000";
		ram_buffer(5855) := X"00000000";
		ram_buffer(5856) := X"00000000";
		ram_buffer(5857) := X"00000000";
		ram_buffer(5858) := X"00000000";
		ram_buffer(5859) := X"00000000";
		ram_buffer(5860) := X"00000000";
		ram_buffer(5861) := X"00000000";
		ram_buffer(5862) := X"00000000";
		ram_buffer(5863) := X"00000000";
		ram_buffer(5864) := X"00000000";
		ram_buffer(5865) := X"00000000";
		ram_buffer(5866) := X"00000000";
		ram_buffer(5867) := X"00000000";
		ram_buffer(5868) := X"00000000";
		ram_buffer(5869) := X"00000000";
		ram_buffer(5870) := X"00000000";
		ram_buffer(5871) := X"00000000";
		ram_buffer(5872) := X"00000000";
		ram_buffer(5873) := X"00000000";
		ram_buffer(5874) := X"00000000";
		ram_buffer(5875) := X"00000000";
		ram_buffer(5876) := X"00000000";
		ram_buffer(5877) := X"00000000";
		ram_buffer(5878) := X"00000000";
		ram_buffer(5879) := X"00000000";
		ram_buffer(5880) := X"00000000";
		ram_buffer(5881) := X"00000000";
		ram_buffer(5882) := X"00000000";
		ram_buffer(5883) := X"00000000";
		ram_buffer(5884) := X"00000000";
		ram_buffer(5885) := X"00000000";
		ram_buffer(5886) := X"00000000";
		ram_buffer(5887) := X"00000000";
		ram_buffer(5888) := X"00000000";
		ram_buffer(5889) := X"00000000";
		ram_buffer(5890) := X"00000000";
		ram_buffer(5891) := X"00000000";
		ram_buffer(5892) := X"00000000";
		ram_buffer(5893) := X"00000000";
		ram_buffer(5894) := X"00000000";
		ram_buffer(5895) := X"00000000";
		ram_buffer(5896) := X"00000000";
		ram_buffer(5897) := X"00000000";
		ram_buffer(5898) := X"00000000";
		ram_buffer(5899) := X"00000000";
		ram_buffer(5900) := X"00000000";
		ram_buffer(5901) := X"00000000";
		ram_buffer(5902) := X"00000000";
		ram_buffer(5903) := X"00000000";
		ram_buffer(5904) := X"00000000";
		ram_buffer(5905) := X"00000000";
		ram_buffer(5906) := X"00000000";
		ram_buffer(5907) := X"00000000";
		ram_buffer(5908) := X"00000000";
		ram_buffer(5909) := X"00000000";
		ram_buffer(5910) := X"00000000";
		ram_buffer(5911) := X"00000000";
		ram_buffer(5912) := X"00000000";
		ram_buffer(5913) := X"00000000";
		ram_buffer(5914) := X"00000000";
		ram_buffer(5915) := X"00000000";
		ram_buffer(5916) := X"00000000";
		ram_buffer(5917) := X"00000000";
		ram_buffer(5918) := X"00000000";
		ram_buffer(5919) := X"00000000";
		ram_buffer(5920) := X"00000000";
		ram_buffer(5921) := X"00000000";
		ram_buffer(5922) := X"00000000";
		ram_buffer(5923) := X"00000000";
		ram_buffer(5924) := X"00000000";
		ram_buffer(5925) := X"00000000";
		ram_buffer(5926) := X"00000000";
		ram_buffer(5927) := X"00000000";
		ram_buffer(5928) := X"00000000";
		ram_buffer(5929) := X"00000000";
		ram_buffer(5930) := X"00000000";
		ram_buffer(5931) := X"00000000";
		ram_buffer(5932) := X"00000000";
		ram_buffer(5933) := X"00000000";
		ram_buffer(5934) := X"00000000";
		ram_buffer(5935) := X"00000000";
		ram_buffer(5936) := X"00000000";
		ram_buffer(5937) := X"00000000";
		ram_buffer(5938) := X"00000000";
		ram_buffer(5939) := X"00000000";
		ram_buffer(5940) := X"00000000";
		ram_buffer(5941) := X"00000000";
		ram_buffer(5942) := X"00000000";
		ram_buffer(5943) := X"00000000";
		ram_buffer(5944) := X"00000000";
		ram_buffer(5945) := X"00000000";
		ram_buffer(5946) := X"00000000";
		ram_buffer(5947) := X"00000000";
		ram_buffer(5948) := X"00000000";
		ram_buffer(5949) := X"00000000";
		ram_buffer(5950) := X"00000000";
		ram_buffer(5951) := X"00000000";
		ram_buffer(5952) := X"00000000";
		ram_buffer(5953) := X"00000000";
		ram_buffer(5954) := X"00000000";
		ram_buffer(5955) := X"00000000";
		ram_buffer(5956) := X"00000000";
		ram_buffer(5957) := X"00000000";
		ram_buffer(5958) := X"00000000";
		ram_buffer(5959) := X"00000000";
		ram_buffer(5960) := X"00000000";
		ram_buffer(5961) := X"00000000";
		ram_buffer(5962) := X"00000000";
		ram_buffer(5963) := X"00000000";
		ram_buffer(5964) := X"00000000";
		ram_buffer(5965) := X"00000000";
		ram_buffer(5966) := X"00000000";
		ram_buffer(5967) := X"00000000";
		ram_buffer(5968) := X"00000000";
		ram_buffer(5969) := X"00000000";
		ram_buffer(5970) := X"00000000";
		ram_buffer(5971) := X"00000000";
		ram_buffer(5972) := X"00000000";
		ram_buffer(5973) := X"00000000";
		ram_buffer(5974) := X"00000000";
		ram_buffer(5975) := X"00000000";
		ram_buffer(5976) := X"00000000";
		ram_buffer(5977) := X"00000000";
		ram_buffer(5978) := X"00000000";
		ram_buffer(5979) := X"00000000";
		ram_buffer(5980) := X"00000000";
		ram_buffer(5981) := X"00000000";
		ram_buffer(5982) := X"00000000";
		ram_buffer(5983) := X"00000000";
		ram_buffer(5984) := X"00000000";
		ram_buffer(5985) := X"00000000";
		ram_buffer(5986) := X"00000000";
		ram_buffer(5987) := X"00000000";
		ram_buffer(5988) := X"00000000";
		ram_buffer(5989) := X"00000000";
		ram_buffer(5990) := X"00000000";
		ram_buffer(5991) := X"00000000";
		ram_buffer(5992) := X"00000000";
		ram_buffer(5993) := X"00000000";
		ram_buffer(5994) := X"00000000";
		ram_buffer(5995) := X"00000000";
		ram_buffer(5996) := X"00000000";
		ram_buffer(5997) := X"00000000";
		ram_buffer(5998) := X"00000000";
		ram_buffer(5999) := X"00000000";
		ram_buffer(6000) := X"00000000";
		ram_buffer(6001) := X"00000000";
		ram_buffer(6002) := X"00000000";
		ram_buffer(6003) := X"00000000";
		ram_buffer(6004) := X"00000000";
		ram_buffer(6005) := X"00000000";
		ram_buffer(6006) := X"00000000";
		ram_buffer(6007) := X"00000000";
		ram_buffer(6008) := X"00000000";
		ram_buffer(6009) := X"00000000";
		ram_buffer(6010) := X"00000000";
		ram_buffer(6011) := X"00000000";
		ram_buffer(6012) := X"00000000";
		ram_buffer(6013) := X"00000000";
		ram_buffer(6014) := X"00000000";
		ram_buffer(6015) := X"00000000";
		ram_buffer(6016) := X"00000000";
		ram_buffer(6017) := X"00000000";
		ram_buffer(6018) := X"00000000";
		ram_buffer(6019) := X"00000000";
		ram_buffer(6020) := X"00000000";
		ram_buffer(6021) := X"00000000";
		ram_buffer(6022) := X"00000000";
		ram_buffer(6023) := X"00000000";
		ram_buffer(6024) := X"00000000";
		ram_buffer(6025) := X"00000000";
		ram_buffer(6026) := X"00000000";
		ram_buffer(6027) := X"00000000";
		ram_buffer(6028) := X"00000000";
		ram_buffer(6029) := X"00000000";
		ram_buffer(6030) := X"00000000";
		ram_buffer(6031) := X"00000000";
		ram_buffer(6032) := X"00000000";
		ram_buffer(6033) := X"00000000";
		ram_buffer(6034) := X"00000000";
		ram_buffer(6035) := X"00000000";
		ram_buffer(6036) := X"00000000";
		ram_buffer(6037) := X"00000000";
		ram_buffer(6038) := X"00000000";
		ram_buffer(6039) := X"00000000";
		ram_buffer(6040) := X"00000000";
		ram_buffer(6041) := X"00000000";
		ram_buffer(6042) := X"00000000";
		ram_buffer(6043) := X"00000000";
		ram_buffer(6044) := X"00000000";
		ram_buffer(6045) := X"00000000";
		ram_buffer(6046) := X"00000000";
		ram_buffer(6047) := X"00000000";
		ram_buffer(6048) := X"00000000";
		ram_buffer(6049) := X"00000000";
		ram_buffer(6050) := X"00000000";
		ram_buffer(6051) := X"00000000";
		ram_buffer(6052) := X"00000000";
		ram_buffer(6053) := X"00000000";
		ram_buffer(6054) := X"00000000";
		ram_buffer(6055) := X"00000000";
		ram_buffer(6056) := X"00000000";
		ram_buffer(6057) := X"00000000";
		ram_buffer(6058) := X"00000000";
		ram_buffer(6059) := X"00000000";
		ram_buffer(6060) := X"00000000";
		ram_buffer(6061) := X"00000000";
		ram_buffer(6062) := X"00000000";
		ram_buffer(6063) := X"00000000";
		ram_buffer(6064) := X"00000000";
		ram_buffer(6065) := X"00000000";
		ram_buffer(6066) := X"00000000";
		ram_buffer(6067) := X"00000000";
		ram_buffer(6068) := X"00000000";
		ram_buffer(6069) := X"00000000";
		ram_buffer(6070) := X"00000000";
		ram_buffer(6071) := X"00000000";
		ram_buffer(6072) := X"00000000";
		ram_buffer(6073) := X"00000000";
		ram_buffer(6074) := X"00000000";
		ram_buffer(6075) := X"00000000";
		ram_buffer(6076) := X"00000000";
		ram_buffer(6077) := X"00000000";
		ram_buffer(6078) := X"00000000";
		ram_buffer(6079) := X"00000000";
		ram_buffer(6080) := X"00000000";
		ram_buffer(6081) := X"00000000";
		ram_buffer(6082) := X"00000000";
		ram_buffer(6083) := X"00000000";
		ram_buffer(6084) := X"00000000";
		ram_buffer(6085) := X"00000000";
		ram_buffer(6086) := X"00000000";
		ram_buffer(6087) := X"00000000";
		ram_buffer(6088) := X"00000000";
		ram_buffer(6089) := X"00000000";
		ram_buffer(6090) := X"00000000";
		ram_buffer(6091) := X"00000000";
		ram_buffer(6092) := X"00000000";
		ram_buffer(6093) := X"00000000";
		ram_buffer(6094) := X"00000000";
		ram_buffer(6095) := X"00000000";
		ram_buffer(6096) := X"00000000";
		ram_buffer(6097) := X"00000000";
		ram_buffer(6098) := X"00000000";
		ram_buffer(6099) := X"00000000";
		ram_buffer(6100) := X"00000000";
		ram_buffer(6101) := X"00000000";
		ram_buffer(6102) := X"00000000";
		ram_buffer(6103) := X"00000000";
		ram_buffer(6104) := X"00000000";
		ram_buffer(6105) := X"00000000";
		ram_buffer(6106) := X"00000000";
		ram_buffer(6107) := X"00000000";
		ram_buffer(6108) := X"00000000";
		ram_buffer(6109) := X"00000000";
		ram_buffer(6110) := X"00000000";
		ram_buffer(6111) := X"00000000";
		ram_buffer(6112) := X"00000000";
		ram_buffer(6113) := X"00000000";
		ram_buffer(6114) := X"00000000";
		ram_buffer(6115) := X"00000000";
		ram_buffer(6116) := X"00000000";
		ram_buffer(6117) := X"00000000";
		ram_buffer(6118) := X"00000000";
		ram_buffer(6119) := X"00000000";
		ram_buffer(6120) := X"00000000";
		ram_buffer(6121) := X"00000000";
		ram_buffer(6122) := X"00000000";
		ram_buffer(6123) := X"00000000";
		ram_buffer(6124) := X"00000000";
		ram_buffer(6125) := X"00000000";
		ram_buffer(6126) := X"00000000";
		ram_buffer(6127) := X"00000000";
		ram_buffer(6128) := X"00000000";
		ram_buffer(6129) := X"00000000";
		ram_buffer(6130) := X"00000000";
		ram_buffer(6131) := X"00000000";
		ram_buffer(6132) := X"00000000";
		ram_buffer(6133) := X"00000000";
		ram_buffer(6134) := X"00000000";
		ram_buffer(6135) := X"00000000";
		ram_buffer(6136) := X"00000000";
		ram_buffer(6137) := X"00000000";
		ram_buffer(6138) := X"00000000";
		ram_buffer(6139) := X"00000000";
		ram_buffer(6140) := X"00000000";
		ram_buffer(6141) := X"00000000";
		ram_buffer(6142) := X"00000000";
		ram_buffer(6143) := X"00000000";
		ram_buffer(6144) := X"00000000";
		ram_buffer(6145) := X"00000000";
		ram_buffer(6146) := X"00000000";
		ram_buffer(6147) := X"00000000";
		ram_buffer(6148) := X"00000000";
		ram_buffer(6149) := X"00000000";
		ram_buffer(6150) := X"00000000";
		ram_buffer(6151) := X"00000000";
		ram_buffer(6152) := X"00000000";
		ram_buffer(6153) := X"00000000";
		ram_buffer(6154) := X"00000000";
		ram_buffer(6155) := X"00000000";
		ram_buffer(6156) := X"00000000";
		ram_buffer(6157) := X"00000000";
		ram_buffer(6158) := X"00000000";
		ram_buffer(6159) := X"00000000";
		ram_buffer(6160) := X"00000000";
		ram_buffer(6161) := X"00000000";
		ram_buffer(6162) := X"00000000";
		ram_buffer(6163) := X"00000000";
		ram_buffer(6164) := X"00000000";
		ram_buffer(6165) := X"00000000";
		ram_buffer(6166) := X"00000000";
		ram_buffer(6167) := X"00000000";
		ram_buffer(6168) := X"00000000";
		ram_buffer(6169) := X"00000000";
		ram_buffer(6170) := X"00000000";
		ram_buffer(6171) := X"00000000";
		ram_buffer(6172) := X"00000000";
		ram_buffer(6173) := X"00000000";
		ram_buffer(6174) := X"00000000";
		ram_buffer(6175) := X"00000000";
		ram_buffer(6176) := X"00000000";
		ram_buffer(6177) := X"00000000";
		ram_buffer(6178) := X"00000000";
		ram_buffer(6179) := X"00000000";
		ram_buffer(6180) := X"00000000";
		ram_buffer(6181) := X"00000000";
		ram_buffer(6182) := X"00000000";
		ram_buffer(6183) := X"00000000";
		ram_buffer(6184) := X"00000000";
		ram_buffer(6185) := X"00000000";
		ram_buffer(6186) := X"00000000";
		ram_buffer(6187) := X"00000000";
		ram_buffer(6188) := X"00000000";
		ram_buffer(6189) := X"00000000";
		ram_buffer(6190) := X"00000000";
		ram_buffer(6191) := X"00000000";
		ram_buffer(6192) := X"00000000";
		ram_buffer(6193) := X"00000000";
		ram_buffer(6194) := X"00000000";
		ram_buffer(6195) := X"00000000";
		ram_buffer(6196) := X"00000000";
		ram_buffer(6197) := X"00000000";
		ram_buffer(6198) := X"00000000";
		ram_buffer(6199) := X"00000000";
		ram_buffer(6200) := X"00000000";
		ram_buffer(6201) := X"00000000";
		ram_buffer(6202) := X"00000000";
		ram_buffer(6203) := X"00000000";
		ram_buffer(6204) := X"00000000";
		ram_buffer(6205) := X"00000000";
		ram_buffer(6206) := X"00000000";
		ram_buffer(6207) := X"00000000";
		ram_buffer(6208) := X"00000000";
		ram_buffer(6209) := X"00000000";
		ram_buffer(6210) := X"00000000";
		ram_buffer(6211) := X"00000000";
		ram_buffer(6212) := X"00000000";
		ram_buffer(6213) := X"00000000";
		ram_buffer(6214) := X"00000000";
		ram_buffer(6215) := X"00000000";
		ram_buffer(6216) := X"00000000";
		ram_buffer(6217) := X"00000000";
		ram_buffer(6218) := X"00000000";
		ram_buffer(6219) := X"00000000";
		ram_buffer(6220) := X"00000000";
		ram_buffer(6221) := X"00000000";
		ram_buffer(6222) := X"00000000";
		ram_buffer(6223) := X"00000000";
		ram_buffer(6224) := X"00000000";
		ram_buffer(6225) := X"00000000";
		ram_buffer(6226) := X"00000000";
		ram_buffer(6227) := X"00000000";
		ram_buffer(6228) := X"00000000";
		ram_buffer(6229) := X"00000000";
		ram_buffer(6230) := X"00000000";
		ram_buffer(6231) := X"00000000";
		ram_buffer(6232) := X"00000000";
		ram_buffer(6233) := X"00000000";
		ram_buffer(6234) := X"00000000";
		ram_buffer(6235) := X"00000000";
		ram_buffer(6236) := X"00000000";
		ram_buffer(6237) := X"00000000";
		ram_buffer(6238) := X"00000000";
		ram_buffer(6239) := X"00000000";
		ram_buffer(6240) := X"00000000";
		ram_buffer(6241) := X"00000000";
		ram_buffer(6242) := X"00000000";
		ram_buffer(6243) := X"00000000";
		ram_buffer(6244) := X"00000000";
		ram_buffer(6245) := X"00000000";
		ram_buffer(6246) := X"00000000";
		ram_buffer(6247) := X"00000000";
		ram_buffer(6248) := X"00000000";
		ram_buffer(6249) := X"00000000";
		ram_buffer(6250) := X"00000000";
		ram_buffer(6251) := X"00000000";
		ram_buffer(6252) := X"00000000";
		ram_buffer(6253) := X"00000000";
		ram_buffer(6254) := X"00000000";
		ram_buffer(6255) := X"00000000";
		ram_buffer(6256) := X"00000000";
		ram_buffer(6257) := X"00000000";
		ram_buffer(6258) := X"00000000";
		ram_buffer(6259) := X"00000000";
		ram_buffer(6260) := X"00000000";
		ram_buffer(6261) := X"00000000";
		ram_buffer(6262) := X"00000000";
		ram_buffer(6263) := X"00000000";
		ram_buffer(6264) := X"00000000";
		ram_buffer(6265) := X"00000000";
		ram_buffer(6266) := X"00000000";
		ram_buffer(6267) := X"00000000";
		ram_buffer(6268) := X"00000000";
		ram_buffer(6269) := X"00000000";
		ram_buffer(6270) := X"00000000";
		ram_buffer(6271) := X"00000000";
		ram_buffer(6272) := X"00000000";
		ram_buffer(6273) := X"00000000";
		ram_buffer(6274) := X"00000000";
		ram_buffer(6275) := X"00000000";
		ram_buffer(6276) := X"00000000";
		ram_buffer(6277) := X"00000000";
		ram_buffer(6278) := X"00000000";
		ram_buffer(6279) := X"00000000";
		ram_buffer(6280) := X"00000000";
		ram_buffer(6281) := X"00000000";
		ram_buffer(6282) := X"00000000";
		ram_buffer(6283) := X"00000000";
		ram_buffer(6284) := X"00000000";
		ram_buffer(6285) := X"00000000";
		ram_buffer(6286) := X"00000000";
		ram_buffer(6287) := X"00000000";
		ram_buffer(6288) := X"00000000";
		ram_buffer(6289) := X"00000000";
		ram_buffer(6290) := X"00000000";
		ram_buffer(6291) := X"00000000";
		ram_buffer(6292) := X"00000000";
		ram_buffer(6293) := X"00000000";
		ram_buffer(6294) := X"00000000";
		ram_buffer(6295) := X"00000000";
		ram_buffer(6296) := X"00000000";
		ram_buffer(6297) := X"00000000";
		ram_buffer(6298) := X"00000000";
		ram_buffer(6299) := X"00000000";
		ram_buffer(6300) := X"00000000";
		ram_buffer(6301) := X"00000000";
		ram_buffer(6302) := X"00000000";
		ram_buffer(6303) := X"00000000";
		ram_buffer(6304) := X"00000000";
		ram_buffer(6305) := X"00000000";
		ram_buffer(6306) := X"00000000";
		ram_buffer(6307) := X"00000000";
		ram_buffer(6308) := X"00000000";
		ram_buffer(6309) := X"00000000";
		ram_buffer(6310) := X"00000000";
		ram_buffer(6311) := X"00000000";
		ram_buffer(6312) := X"00000000";
		ram_buffer(6313) := X"00000000";
		ram_buffer(6314) := X"00000000";
		ram_buffer(6315) := X"00000000";
		ram_buffer(6316) := X"00000000";
		ram_buffer(6317) := X"00000000";
		ram_buffer(6318) := X"00000000";
		ram_buffer(6319) := X"00000000";
		ram_buffer(6320) := X"00000000";
		ram_buffer(6321) := X"00000000";
		ram_buffer(6322) := X"00000000";
		ram_buffer(6323) := X"00000000";
		ram_buffer(6324) := X"00000000";
		ram_buffer(6325) := X"00000000";
		ram_buffer(6326) := X"00000000";
		ram_buffer(6327) := X"00000000";
		ram_buffer(6328) := X"00000000";
		ram_buffer(6329) := X"00000000";
		ram_buffer(6330) := X"00000000";
		ram_buffer(6331) := X"00000000";
		ram_buffer(6332) := X"00000000";
		ram_buffer(6333) := X"00000000";
		ram_buffer(6334) := X"00000000";
		ram_buffer(6335) := X"00000000";
		ram_buffer(6336) := X"00000000";
		ram_buffer(6337) := X"00000000";
		ram_buffer(6338) := X"00000000";
		ram_buffer(6339) := X"00000000";
		ram_buffer(6340) := X"00000000";
		ram_buffer(6341) := X"00000000";
		ram_buffer(6342) := X"00000000";
		ram_buffer(6343) := X"00000000";
		ram_buffer(6344) := X"00000000";
		ram_buffer(6345) := X"00000000";
		ram_buffer(6346) := X"00000000";
		ram_buffer(6347) := X"00000000";
		ram_buffer(6348) := X"00000000";
		ram_buffer(6349) := X"00000000";
		ram_buffer(6350) := X"00000000";
		ram_buffer(6351) := X"00000000";
		ram_buffer(6352) := X"00000000";
		ram_buffer(6353) := X"00000000";
		ram_buffer(6354) := X"00000000";
		ram_buffer(6355) := X"00000000";
		ram_buffer(6356) := X"00000000";
		ram_buffer(6357) := X"00000000";
		ram_buffer(6358) := X"00000000";
		ram_buffer(6359) := X"00000000";
		ram_buffer(6360) := X"00000000";
		ram_buffer(6361) := X"00000000";
		ram_buffer(6362) := X"00000000";
		ram_buffer(6363) := X"00000000";
		ram_buffer(6364) := X"00000000";
		ram_buffer(6365) := X"00000000";
		ram_buffer(6366) := X"00000000";
		ram_buffer(6367) := X"00000000";
		ram_buffer(6368) := X"00000000";
		ram_buffer(6369) := X"00000000";
		ram_buffer(6370) := X"00000000";
		ram_buffer(6371) := X"00000000";
		ram_buffer(6372) := X"00000000";
		ram_buffer(6373) := X"00000000";
		ram_buffer(6374) := X"00000000";
		ram_buffer(6375) := X"00000000";
		ram_buffer(6376) := X"00000000";
		ram_buffer(6377) := X"00000000";
		ram_buffer(6378) := X"00000000";
		ram_buffer(6379) := X"00000000";
		ram_buffer(6380) := X"00000000";
		ram_buffer(6381) := X"00000000";
		ram_buffer(6382) := X"00000000";
		ram_buffer(6383) := X"00000000";
		ram_buffer(6384) := X"00000000";
		ram_buffer(6385) := X"00000000";
		ram_buffer(6386) := X"00000000";
		ram_buffer(6387) := X"00000000";
		ram_buffer(6388) := X"00000000";
		ram_buffer(6389) := X"00000000";
		ram_buffer(6390) := X"00000000";
		ram_buffer(6391) := X"00000000";
		ram_buffer(6392) := X"00000000";
		ram_buffer(6393) := X"00000000";
		ram_buffer(6394) := X"00000000";
		ram_buffer(6395) := X"00000000";
		ram_buffer(6396) := X"00000000";
		ram_buffer(6397) := X"00000000";
		ram_buffer(6398) := X"00000000";
		ram_buffer(6399) := X"00000000";
		ram_buffer(6400) := X"00000000";
		ram_buffer(6401) := X"00000000";
		ram_buffer(6402) := X"00000000";
		ram_buffer(6403) := X"00000000";
		ram_buffer(6404) := X"00000000";
		ram_buffer(6405) := X"00000000";
		ram_buffer(6406) := X"00000000";
		ram_buffer(6407) := X"00000000";
		ram_buffer(6408) := X"00000000";
		ram_buffer(6409) := X"00000000";
		ram_buffer(6410) := X"00000000";
		ram_buffer(6411) := X"00000000";
		ram_buffer(6412) := X"00000000";
		ram_buffer(6413) := X"00000000";
		ram_buffer(6414) := X"00000000";
		ram_buffer(6415) := X"00000000";
		ram_buffer(6416) := X"00000000";
		ram_buffer(6417) := X"00000000";
		ram_buffer(6418) := X"00000000";
		ram_buffer(6419) := X"00000000";
		ram_buffer(6420) := X"00000000";
		ram_buffer(6421) := X"00000000";
		ram_buffer(6422) := X"00000000";
		ram_buffer(6423) := X"00000000";
		ram_buffer(6424) := X"00000000";
		ram_buffer(6425) := X"00000000";
		ram_buffer(6426) := X"00000000";
		ram_buffer(6427) := X"00000000";
		ram_buffer(6428) := X"00000000";
		ram_buffer(6429) := X"00000000";
		ram_buffer(6430) := X"00000000";
		ram_buffer(6431) := X"00000000";
		ram_buffer(6432) := X"00000000";
		ram_buffer(6433) := X"00000000";
		ram_buffer(6434) := X"00000000";
		ram_buffer(6435) := X"00000000";
		ram_buffer(6436) := X"00000000";
		ram_buffer(6437) := X"00000000";
		ram_buffer(6438) := X"00000000";
		ram_buffer(6439) := X"00000000";
		ram_buffer(6440) := X"00000000";
		ram_buffer(6441) := X"00000000";
		ram_buffer(6442) := X"00000000";
		ram_buffer(6443) := X"00000000";
		ram_buffer(6444) := X"00000000";
		ram_buffer(6445) := X"00000000";
		ram_buffer(6446) := X"00000000";
		ram_buffer(6447) := X"00000000";
		ram_buffer(6448) := X"00000000";
		ram_buffer(6449) := X"00000000";
		ram_buffer(6450) := X"00000000";
		ram_buffer(6451) := X"00000000";
		ram_buffer(6452) := X"00000000";
		ram_buffer(6453) := X"00000000";
		ram_buffer(6454) := X"00000000";
		ram_buffer(6455) := X"00000000";
		ram_buffer(6456) := X"00000000";
		ram_buffer(6457) := X"00000000";
		ram_buffer(6458) := X"00000000";
		ram_buffer(6459) := X"00000000";
		ram_buffer(6460) := X"00000000";
		ram_buffer(6461) := X"00000000";
		ram_buffer(6462) := X"00000000";
		ram_buffer(6463) := X"00000000";
		ram_buffer(6464) := X"00000000";
		ram_buffer(6465) := X"00000000";
		ram_buffer(6466) := X"00000000";
		ram_buffer(6467) := X"00000000";
		ram_buffer(6468) := X"00000000";
		ram_buffer(6469) := X"00000000";
		ram_buffer(6470) := X"00000000";
		ram_buffer(6471) := X"00000000";
		ram_buffer(6472) := X"00000000";
		ram_buffer(6473) := X"00000000";
		ram_buffer(6474) := X"00000000";
		ram_buffer(6475) := X"00000000";
		ram_buffer(6476) := X"00000000";
		ram_buffer(6477) := X"00000000";
		ram_buffer(6478) := X"00000000";
		ram_buffer(6479) := X"00000000";
		ram_buffer(6480) := X"00000000";
		ram_buffer(6481) := X"00000000";
		ram_buffer(6482) := X"00000000";
		ram_buffer(6483) := X"00000000";
		ram_buffer(6484) := X"00000000";
		ram_buffer(6485) := X"00000000";
		ram_buffer(6486) := X"00000000";
		ram_buffer(6487) := X"00000000";
		ram_buffer(6488) := X"00000000";
		ram_buffer(6489) := X"00000000";
		ram_buffer(6490) := X"00000000";
		ram_buffer(6491) := X"00000000";
		ram_buffer(6492) := X"00000000";
		ram_buffer(6493) := X"00000000";
		ram_buffer(6494) := X"00000000";
		ram_buffer(6495) := X"00000000";
		ram_buffer(6496) := X"00000000";
		ram_buffer(6497) := X"00000000";
		ram_buffer(6498) := X"00000000";
		ram_buffer(6499) := X"00000000";
		ram_buffer(6500) := X"00000000";
		ram_buffer(6501) := X"00000000";
		ram_buffer(6502) := X"00000000";
		ram_buffer(6503) := X"00000000";
		ram_buffer(6504) := X"00000000";
		ram_buffer(6505) := X"00000000";
		ram_buffer(6506) := X"00000000";
		ram_buffer(6507) := X"00000000";
		ram_buffer(6508) := X"00000000";
		ram_buffer(6509) := X"00000000";
		ram_buffer(6510) := X"00000000";
		ram_buffer(6511) := X"00000000";
		ram_buffer(6512) := X"00000000";
		ram_buffer(6513) := X"00000000";
		ram_buffer(6514) := X"00000000";
		ram_buffer(6515) := X"00000000";
		ram_buffer(6516) := X"00000000";
		ram_buffer(6517) := X"00000000";
		ram_buffer(6518) := X"00000000";
		ram_buffer(6519) := X"00000000";
		ram_buffer(6520) := X"00000000";
		ram_buffer(6521) := X"00000000";
		ram_buffer(6522) := X"00000000";
		ram_buffer(6523) := X"00000000";
		ram_buffer(6524) := X"00000000";
		ram_buffer(6525) := X"00000000";
		ram_buffer(6526) := X"00000000";
		ram_buffer(6527) := X"00000000";
		ram_buffer(6528) := X"00000000";
		ram_buffer(6529) := X"00000000";
		ram_buffer(6530) := X"00000000";
		ram_buffer(6531) := X"00000000";
		ram_buffer(6532) := X"00000000";
		ram_buffer(6533) := X"00000000";
		ram_buffer(6534) := X"00000000";
		ram_buffer(6535) := X"00000000";
		ram_buffer(6536) := X"00000000";
		ram_buffer(6537) := X"00000000";
		ram_buffer(6538) := X"00000000";
		ram_buffer(6539) := X"00000000";
		ram_buffer(6540) := X"00000000";
		ram_buffer(6541) := X"00000000";
		ram_buffer(6542) := X"00000000";
		ram_buffer(6543) := X"00000000";
		ram_buffer(6544) := X"00000000";
		ram_buffer(6545) := X"00000000";
		ram_buffer(6546) := X"00000000";
		ram_buffer(6547) := X"00000000";
		ram_buffer(6548) := X"00000000";
		ram_buffer(6549) := X"00000000";
		ram_buffer(6550) := X"00000000";
		ram_buffer(6551) := X"00000000";
		ram_buffer(6552) := X"00000000";
		ram_buffer(6553) := X"00000000";
		ram_buffer(6554) := X"00000000";
		ram_buffer(6555) := X"00000000";
		ram_buffer(6556) := X"00000000";
		ram_buffer(6557) := X"00000000";
		ram_buffer(6558) := X"00000000";
		ram_buffer(6559) := X"00000000";
		ram_buffer(6560) := X"00000000";
		ram_buffer(6561) := X"00000000";
		ram_buffer(6562) := X"00000000";
		ram_buffer(6563) := X"00000000";
		ram_buffer(6564) := X"00000000";
		ram_buffer(6565) := X"00000000";
		ram_buffer(6566) := X"00000000";
		ram_buffer(6567) := X"00000000";
		ram_buffer(6568) := X"00000000";
		ram_buffer(6569) := X"00000000";
		ram_buffer(6570) := X"00000000";
		ram_buffer(6571) := X"00000000";
		ram_buffer(6572) := X"00000000";
		ram_buffer(6573) := X"00000000";
		ram_buffer(6574) := X"00000000";
		ram_buffer(6575) := X"00000000";
		ram_buffer(6576) := X"00000000";
		ram_buffer(6577) := X"00000000";
		ram_buffer(6578) := X"00000000";
		ram_buffer(6579) := X"00000000";
		ram_buffer(6580) := X"00000000";
		ram_buffer(6581) := X"00000000";
		ram_buffer(6582) := X"00000000";
		ram_buffer(6583) := X"00000000";
		ram_buffer(6584) := X"00000000";
		ram_buffer(6585) := X"00000000";
		ram_buffer(6586) := X"00000000";
		ram_buffer(6587) := X"00000000";
		ram_buffer(6588) := X"00000000";
		ram_buffer(6589) := X"00000000";
		ram_buffer(6590) := X"00000000";
		ram_buffer(6591) := X"00000000";
		ram_buffer(6592) := X"00000000";
		ram_buffer(6593) := X"00000000";
		ram_buffer(6594) := X"00000000";
		ram_buffer(6595) := X"00000000";
		ram_buffer(6596) := X"00000000";
		ram_buffer(6597) := X"00000000";
		ram_buffer(6598) := X"00000000";
		ram_buffer(6599) := X"00000000";
		ram_buffer(6600) := X"00000000";
		ram_buffer(6601) := X"00000000";
		ram_buffer(6602) := X"00000000";
		ram_buffer(6603) := X"00000000";
		ram_buffer(6604) := X"00000000";
		ram_buffer(6605) := X"00000000";
		ram_buffer(6606) := X"00000000";
		ram_buffer(6607) := X"00000000";
		ram_buffer(6608) := X"00000000";
		ram_buffer(6609) := X"00000000";
		ram_buffer(6610) := X"00000000";
		ram_buffer(6611) := X"00000000";
		ram_buffer(6612) := X"00000000";
		ram_buffer(6613) := X"00000000";
		ram_buffer(6614) := X"00000000";
		ram_buffer(6615) := X"00000000";
		ram_buffer(6616) := X"00000000";
		ram_buffer(6617) := X"00000000";
		ram_buffer(6618) := X"00000000";
		ram_buffer(6619) := X"00000000";
		ram_buffer(6620) := X"00000000";
		ram_buffer(6621) := X"00000000";
		ram_buffer(6622) := X"00000000";
		ram_buffer(6623) := X"00000000";
		ram_buffer(6624) := X"00000000";
		ram_buffer(6625) := X"00000000";
		ram_buffer(6626) := X"00000000";
		ram_buffer(6627) := X"00000000";
		ram_buffer(6628) := X"00000000";
		ram_buffer(6629) := X"00000000";
		ram_buffer(6630) := X"00000000";
		ram_buffer(6631) := X"00000000";
		ram_buffer(6632) := X"00000000";
		ram_buffer(6633) := X"00000000";
		ram_buffer(6634) := X"00000000";
		ram_buffer(6635) := X"00000000";
		ram_buffer(6636) := X"00000000";
		ram_buffer(6637) := X"00000000";
		ram_buffer(6638) := X"00000000";
		ram_buffer(6639) := X"00000000";
		ram_buffer(6640) := X"00000000";
		ram_buffer(6641) := X"00000000";
		ram_buffer(6642) := X"00000000";
		ram_buffer(6643) := X"00000000";
		ram_buffer(6644) := X"00000000";
		ram_buffer(6645) := X"00000000";
		ram_buffer(6646) := X"00000000";
		ram_buffer(6647) := X"00000000";
		ram_buffer(6648) := X"00000000";
		ram_buffer(6649) := X"00000000";
		ram_buffer(6650) := X"00000000";
		ram_buffer(6651) := X"00000000";
		ram_buffer(6652) := X"00000000";
		ram_buffer(6653) := X"00000000";
		ram_buffer(6654) := X"00000000";
		ram_buffer(6655) := X"00000000";
		ram_buffer(6656) := X"00000000";
		ram_buffer(6657) := X"00000000";
		ram_buffer(6658) := X"00000000";
		ram_buffer(6659) := X"00000000";
		ram_buffer(6660) := X"00000000";
		ram_buffer(6661) := X"00000000";
		ram_buffer(6662) := X"00000000";
		ram_buffer(6663) := X"00000000";
		ram_buffer(6664) := X"00000000";
		ram_buffer(6665) := X"00000000";
		ram_buffer(6666) := X"00000000";
		ram_buffer(6667) := X"00000000";
		ram_buffer(6668) := X"00000000";
		ram_buffer(6669) := X"00000000";
		ram_buffer(6670) := X"00000000";
		ram_buffer(6671) := X"00000000";
		ram_buffer(6672) := X"00000000";
		ram_buffer(6673) := X"00000000";
		ram_buffer(6674) := X"00000000";
		ram_buffer(6675) := X"00000000";
		ram_buffer(6676) := X"00000000";
		ram_buffer(6677) := X"00000000";
		ram_buffer(6678) := X"00000000";
		ram_buffer(6679) := X"00000000";
		ram_buffer(6680) := X"00000000";
		ram_buffer(6681) := X"00000000";
		ram_buffer(6682) := X"00000000";
		ram_buffer(6683) := X"00000000";
		ram_buffer(6684) := X"00000000";
		ram_buffer(6685) := X"00000000";
		ram_buffer(6686) := X"00000000";
		ram_buffer(6687) := X"00000000";
		ram_buffer(6688) := X"00000000";
		ram_buffer(6689) := X"00000000";
		ram_buffer(6690) := X"00000000";
		ram_buffer(6691) := X"00000000";
		ram_buffer(6692) := X"00000000";
		ram_buffer(6693) := X"00000000";
		ram_buffer(6694) := X"00000000";
		ram_buffer(6695) := X"00000000";
		ram_buffer(6696) := X"00000000";
		ram_buffer(6697) := X"00000000";
		ram_buffer(6698) := X"00000000";
		ram_buffer(6699) := X"00000000";
		ram_buffer(6700) := X"00000000";
		ram_buffer(6701) := X"00000000";
		ram_buffer(6702) := X"00000000";
		ram_buffer(6703) := X"00000000";
		ram_buffer(6704) := X"00000000";
		ram_buffer(6705) := X"00000000";
		ram_buffer(6706) := X"00000000";
		ram_buffer(6707) := X"00000000";
		ram_buffer(6708) := X"00000000";
		ram_buffer(6709) := X"00000000";
		ram_buffer(6710) := X"00000000";
		ram_buffer(6711) := X"00000000";
		ram_buffer(6712) := X"00000000";
		ram_buffer(6713) := X"00000000";
		ram_buffer(6714) := X"00000000";
		ram_buffer(6715) := X"00000000";
		ram_buffer(6716) := X"00000000";
		ram_buffer(6717) := X"00000000";
		ram_buffer(6718) := X"00000000";
		ram_buffer(6719) := X"00000000";
		ram_buffer(6720) := X"00000000";
		ram_buffer(6721) := X"00000000";
		ram_buffer(6722) := X"00000000";
		ram_buffer(6723) := X"00000000";
		ram_buffer(6724) := X"00000000";
		ram_buffer(6725) := X"00000000";
		ram_buffer(6726) := X"00000000";
		ram_buffer(6727) := X"00000000";
		ram_buffer(6728) := X"00000000";
		ram_buffer(6729) := X"00000000";
		ram_buffer(6730) := X"00000000";
		ram_buffer(6731) := X"00000000";
		ram_buffer(6732) := X"00000000";
		ram_buffer(6733) := X"00000000";
		ram_buffer(6734) := X"00000000";
		ram_buffer(6735) := X"00000000";
		ram_buffer(6736) := X"00000000";
		ram_buffer(6737) := X"00000000";
		ram_buffer(6738) := X"00000000";
		ram_buffer(6739) := X"00000000";
		ram_buffer(6740) := X"00000000";
		ram_buffer(6741) := X"00000000";
		ram_buffer(6742) := X"00000000";
		ram_buffer(6743) := X"00000000";
		ram_buffer(6744) := X"00000000";
		ram_buffer(6745) := X"00000000";
		ram_buffer(6746) := X"00000000";
		ram_buffer(6747) := X"00000000";
		ram_buffer(6748) := X"00000000";
		ram_buffer(6749) := X"00000000";
		ram_buffer(6750) := X"00000000";
		ram_buffer(6751) := X"00000000";
		ram_buffer(6752) := X"00000000";
		ram_buffer(6753) := X"00000000";
		ram_buffer(6754) := X"00000000";
		ram_buffer(6755) := X"00000000";
		ram_buffer(6756) := X"00000000";
		ram_buffer(6757) := X"00000000";
		ram_buffer(6758) := X"00000000";
		ram_buffer(6759) := X"00000000";
		ram_buffer(6760) := X"00000000";
		ram_buffer(6761) := X"00000000";
		ram_buffer(6762) := X"00000000";
		ram_buffer(6763) := X"00000000";
		ram_buffer(6764) := X"00000000";
		ram_buffer(6765) := X"00000000";
		ram_buffer(6766) := X"00000000";
		ram_buffer(6767) := X"00000000";
		ram_buffer(6768) := X"00000000";
		ram_buffer(6769) := X"00000000";
		ram_buffer(6770) := X"00000000";
		ram_buffer(6771) := X"00000000";
		ram_buffer(6772) := X"00000000";
		ram_buffer(6773) := X"00000000";
		ram_buffer(6774) := X"00000000";
		ram_buffer(6775) := X"00000000";
		ram_buffer(6776) := X"00000000";
		ram_buffer(6777) := X"00000000";
		ram_buffer(6778) := X"00000000";
		ram_buffer(6779) := X"00000000";
		ram_buffer(6780) := X"00000000";
		ram_buffer(6781) := X"00000000";
		ram_buffer(6782) := X"00000000";
		ram_buffer(6783) := X"00000000";
		ram_buffer(6784) := X"00000000";
		ram_buffer(6785) := X"00000000";
		ram_buffer(6786) := X"00000000";
		ram_buffer(6787) := X"00000000";
		ram_buffer(6788) := X"00000000";
		ram_buffer(6789) := X"00000000";
		ram_buffer(6790) := X"00000000";
		ram_buffer(6791) := X"00000000";
		ram_buffer(6792) := X"00000000";
		ram_buffer(6793) := X"00000000";
		ram_buffer(6794) := X"00000000";
		ram_buffer(6795) := X"00000000";
		ram_buffer(6796) := X"00000000";
		ram_buffer(6797) := X"00000000";
		ram_buffer(6798) := X"00000000";
		ram_buffer(6799) := X"00000000";
		ram_buffer(6800) := X"00000000";
		ram_buffer(6801) := X"00000000";
		ram_buffer(6802) := X"00000000";
		ram_buffer(6803) := X"00000000";
		ram_buffer(6804) := X"00000000";
		ram_buffer(6805) := X"00000000";
		ram_buffer(6806) := X"00000000";
		ram_buffer(6807) := X"00000000";
		ram_buffer(6808) := X"00000000";
		ram_buffer(6809) := X"00000000";
		ram_buffer(6810) := X"00000000";
		ram_buffer(6811) := X"00000000";
		ram_buffer(6812) := X"00000000";
		ram_buffer(6813) := X"00000000";
		ram_buffer(6814) := X"00000000";
		ram_buffer(6815) := X"00000000";
		ram_buffer(6816) := X"00000000";
		ram_buffer(6817) := X"00000000";
		ram_buffer(6818) := X"00000000";
		ram_buffer(6819) := X"00000000";
		ram_buffer(6820) := X"00000000";
		ram_buffer(6821) := X"00000000";
		ram_buffer(6822) := X"00000000";
		ram_buffer(6823) := X"00000000";
		ram_buffer(6824) := X"00000000";
		ram_buffer(6825) := X"00000000";
		ram_buffer(6826) := X"00000000";
		ram_buffer(6827) := X"00000000";
		ram_buffer(6828) := X"00000000";
		ram_buffer(6829) := X"00000000";
		ram_buffer(6830) := X"00000000";
		ram_buffer(6831) := X"00000000";
		ram_buffer(6832) := X"00000000";
		ram_buffer(6833) := X"00000000";
		ram_buffer(6834) := X"00000000";
		ram_buffer(6835) := X"00000000";
		ram_buffer(6836) := X"00000000";
		ram_buffer(6837) := X"00000000";
		ram_buffer(6838) := X"00000000";
		ram_buffer(6839) := X"00000000";
		ram_buffer(6840) := X"00000000";
		ram_buffer(6841) := X"00000000";
		ram_buffer(6842) := X"00000000";
		ram_buffer(6843) := X"00000000";
		ram_buffer(6844) := X"00000000";
		ram_buffer(6845) := X"00000000";
		ram_buffer(6846) := X"00000000";
		ram_buffer(6847) := X"00000000";
		ram_buffer(6848) := X"00000000";
		ram_buffer(6849) := X"00000000";
		ram_buffer(6850) := X"00000000";
		ram_buffer(6851) := X"00000000";
		ram_buffer(6852) := X"00000000";
		ram_buffer(6853) := X"00000000";
		ram_buffer(6854) := X"00000000";
		ram_buffer(6855) := X"00000000";
		ram_buffer(6856) := X"00000000";
		ram_buffer(6857) := X"00000000";
		ram_buffer(6858) := X"00000000";
		ram_buffer(6859) := X"00000000";
		ram_buffer(6860) := X"00000000";
		ram_buffer(6861) := X"00000000";
		ram_buffer(6862) := X"00000000";
		ram_buffer(6863) := X"00000000";
		ram_buffer(6864) := X"00000000";
		ram_buffer(6865) := X"00000000";
		ram_buffer(6866) := X"00000000";
		ram_buffer(6867) := X"00000000";
		ram_buffer(6868) := X"00000000";
		ram_buffer(6869) := X"00000000";
		ram_buffer(6870) := X"00000000";
		ram_buffer(6871) := X"00000000";
		ram_buffer(6872) := X"00000000";
		ram_buffer(6873) := X"00000000";
		ram_buffer(6874) := X"00000000";
		ram_buffer(6875) := X"00000000";
		ram_buffer(6876) := X"00000000";
		ram_buffer(6877) := X"00000000";
		ram_buffer(6878) := X"00000000";
		ram_buffer(6879) := X"00000000";
		ram_buffer(6880) := X"00000000";
		ram_buffer(6881) := X"00000000";
		ram_buffer(6882) := X"00000000";
		ram_buffer(6883) := X"00000000";
		ram_buffer(6884) := X"00000000";
		ram_buffer(6885) := X"00000000";
		ram_buffer(6886) := X"00000000";
		ram_buffer(6887) := X"00000000";
		ram_buffer(6888) := X"00000000";
		ram_buffer(6889) := X"00000000";
		ram_buffer(6890) := X"00000000";
		ram_buffer(6891) := X"00000000";
		ram_buffer(6892) := X"00000000";
		ram_buffer(6893) := X"00000000";
		ram_buffer(6894) := X"00000000";
		ram_buffer(6895) := X"00000000";
		ram_buffer(6896) := X"00000000";
		ram_buffer(6897) := X"00000000";
		ram_buffer(6898) := X"00000000";
		ram_buffer(6899) := X"00000000";
		ram_buffer(6900) := X"00000000";
		ram_buffer(6901) := X"00000000";
		ram_buffer(6902) := X"00000000";
		ram_buffer(6903) := X"00000000";
		ram_buffer(6904) := X"00000000";
		ram_buffer(6905) := X"00000000";
		ram_buffer(6906) := X"00000000";
		ram_buffer(6907) := X"00000000";
		ram_buffer(6908) := X"00000000";
		ram_buffer(6909) := X"00000000";
		ram_buffer(6910) := X"00000000";
		ram_buffer(6911) := X"00000000";
		ram_buffer(6912) := X"00000000";
		ram_buffer(6913) := X"00000000";
		ram_buffer(6914) := X"00000000";
		ram_buffer(6915) := X"00000000";
		ram_buffer(6916) := X"00000000";
		ram_buffer(6917) := X"00000000";
		ram_buffer(6918) := X"00000000";
		ram_buffer(6919) := X"00000000";
		ram_buffer(6920) := X"00000000";
		ram_buffer(6921) := X"00000000";
		ram_buffer(6922) := X"00000000";
		ram_buffer(6923) := X"00000000";
		ram_buffer(6924) := X"00000000";
		ram_buffer(6925) := X"00000000";
		ram_buffer(6926) := X"00000000";
		ram_buffer(6927) := X"00000000";
		ram_buffer(6928) := X"00000000";
		ram_buffer(6929) := X"00000000";
		ram_buffer(6930) := X"00000000";
		ram_buffer(6931) := X"00000000";
		ram_buffer(6932) := X"00000000";
		ram_buffer(6933) := X"00000000";
		ram_buffer(6934) := X"00000000";
		ram_buffer(6935) := X"00000000";
		ram_buffer(6936) := X"00000000";
		ram_buffer(6937) := X"00000000";
		ram_buffer(6938) := X"00000000";
		ram_buffer(6939) := X"00000000";
		ram_buffer(6940) := X"00000000";
		ram_buffer(6941) := X"00000000";
		ram_buffer(6942) := X"00000000";
		ram_buffer(6943) := X"00000000";
		ram_buffer(6944) := X"00000000";
		ram_buffer(6945) := X"00000000";
		ram_buffer(6946) := X"00000000";
		ram_buffer(6947) := X"00000000";
		ram_buffer(6948) := X"00000000";
		ram_buffer(6949) := X"00000000";
		ram_buffer(6950) := X"00000000";
		ram_buffer(6951) := X"00000000";
		ram_buffer(6952) := X"00000000";
		ram_buffer(6953) := X"00000000";
		ram_buffer(6954) := X"00000000";
		ram_buffer(6955) := X"00000000";
		ram_buffer(6956) := X"00000000";
		ram_buffer(6957) := X"00000000";
		ram_buffer(6958) := X"00000000";
		ram_buffer(6959) := X"00000000";
		ram_buffer(6960) := X"00000000";
		ram_buffer(6961) := X"00000000";
		ram_buffer(6962) := X"00000000";
		ram_buffer(6963) := X"00000000";
		ram_buffer(6964) := X"00000000";
		ram_buffer(6965) := X"00000000";
		ram_buffer(6966) := X"00000000";
		ram_buffer(6967) := X"00000000";
		ram_buffer(6968) := X"00000000";
		ram_buffer(6969) := X"00000000";
		ram_buffer(6970) := X"00000000";
		ram_buffer(6971) := X"00000000";
		ram_buffer(6972) := X"00000000";
		ram_buffer(6973) := X"00000000";
		ram_buffer(6974) := X"00000000";
		ram_buffer(6975) := X"00000000";
		ram_buffer(6976) := X"00000000";
		ram_buffer(6977) := X"00000000";
		ram_buffer(6978) := X"00000000";
		ram_buffer(6979) := X"00000000";
		ram_buffer(6980) := X"00000000";
		ram_buffer(6981) := X"00000000";
		ram_buffer(6982) := X"00000000";
		ram_buffer(6983) := X"00000000";
		ram_buffer(6984) := X"00000000";
		ram_buffer(6985) := X"00000000";
		ram_buffer(6986) := X"00000000";
		ram_buffer(6987) := X"00000000";
		ram_buffer(6988) := X"00000000";
		ram_buffer(6989) := X"00000000";
		ram_buffer(6990) := X"00000000";
		ram_buffer(6991) := X"00000000";
		ram_buffer(6992) := X"00000000";
		ram_buffer(6993) := X"00000000";
		ram_buffer(6994) := X"00000000";
		ram_buffer(6995) := X"00000000";
		ram_buffer(6996) := X"00000000";
		ram_buffer(6997) := X"00000000";
		ram_buffer(6998) := X"00000000";
		ram_buffer(6999) := X"00000000";
		ram_buffer(7000) := X"00000000";
		ram_buffer(7001) := X"00000000";
		ram_buffer(7002) := X"00000000";
		ram_buffer(7003) := X"00000000";
		ram_buffer(7004) := X"00000000";
		ram_buffer(7005) := X"00000000";
		ram_buffer(7006) := X"00000000";
		ram_buffer(7007) := X"00000000";
		ram_buffer(7008) := X"00000000";
		ram_buffer(7009) := X"00000000";
		ram_buffer(7010) := X"00000000";
		ram_buffer(7011) := X"00000000";
		ram_buffer(7012) := X"00000000";
		ram_buffer(7013) := X"00000000";
		ram_buffer(7014) := X"00000000";
		ram_buffer(7015) := X"00000000";
		ram_buffer(7016) := X"00000000";
		ram_buffer(7017) := X"00000000";
		ram_buffer(7018) := X"00000000";
		ram_buffer(7019) := X"00000000";
		ram_buffer(7020) := X"00000000";
		ram_buffer(7021) := X"00000000";
		ram_buffer(7022) := X"00000000";
		ram_buffer(7023) := X"00000000";
		ram_buffer(7024) := X"00000000";
		ram_buffer(7025) := X"00000000";
		ram_buffer(7026) := X"00000000";
		ram_buffer(7027) := X"00000000";
		ram_buffer(7028) := X"00000000";
		ram_buffer(7029) := X"00000000";
		ram_buffer(7030) := X"00000000";
		ram_buffer(7031) := X"00000000";
		ram_buffer(7032) := X"00000000";
		ram_buffer(7033) := X"00000000";
		ram_buffer(7034) := X"00000000";
		ram_buffer(7035) := X"00000000";
		ram_buffer(7036) := X"00000000";
		ram_buffer(7037) := X"00000000";
		ram_buffer(7038) := X"00000000";
		ram_buffer(7039) := X"00000000";
		ram_buffer(7040) := X"00000000";
		ram_buffer(7041) := X"00000000";
		ram_buffer(7042) := X"00000000";
		ram_buffer(7043) := X"00000000";
		ram_buffer(7044) := X"00000000";
		ram_buffer(7045) := X"00000000";
		ram_buffer(7046) := X"00000000";
		ram_buffer(7047) := X"00000000";
		ram_buffer(7048) := X"00000000";
		ram_buffer(7049) := X"00000000";
		ram_buffer(7050) := X"00000000";
		ram_buffer(7051) := X"00000000";
		ram_buffer(7052) := X"00000000";
		ram_buffer(7053) := X"00000000";
		ram_buffer(7054) := X"00000000";
		ram_buffer(7055) := X"00000000";
		ram_buffer(7056) := X"00000000";
		ram_buffer(7057) := X"00000000";
		ram_buffer(7058) := X"00000000";
		ram_buffer(7059) := X"00000000";
		ram_buffer(7060) := X"00000000";
		ram_buffer(7061) := X"00000000";
		ram_buffer(7062) := X"00000000";
		ram_buffer(7063) := X"00000000";
		ram_buffer(7064) := X"00000000";
		ram_buffer(7065) := X"00000000";
		ram_buffer(7066) := X"00000000";
		ram_buffer(7067) := X"00000000";
		ram_buffer(7068) := X"00000000";
		ram_buffer(7069) := X"00000000";
		ram_buffer(7070) := X"00000000";
		ram_buffer(7071) := X"00000000";
		ram_buffer(7072) := X"00000000";
		ram_buffer(7073) := X"00000000";
		ram_buffer(7074) := X"00000000";
		ram_buffer(7075) := X"00000000";
		ram_buffer(7076) := X"00000000";
		ram_buffer(7077) := X"00000000";
		ram_buffer(7078) := X"00000000";
		ram_buffer(7079) := X"00000000";
		ram_buffer(7080) := X"00000000";
		ram_buffer(7081) := X"00000000";
		ram_buffer(7082) := X"00000000";
		ram_buffer(7083) := X"00000000";
		ram_buffer(7084) := X"00000000";
		ram_buffer(7085) := X"00000000";
		ram_buffer(7086) := X"00000000";
		ram_buffer(7087) := X"00000000";
		ram_buffer(7088) := X"00000000";
		ram_buffer(7089) := X"00000000";
		ram_buffer(7090) := X"00000000";
		ram_buffer(7091) := X"00000000";
		ram_buffer(7092) := X"00000000";
		ram_buffer(7093) := X"00000000";
		ram_buffer(7094) := X"00000000";
		ram_buffer(7095) := X"00000000";
		ram_buffer(7096) := X"00000000";
		ram_buffer(7097) := X"00000000";
		ram_buffer(7098) := X"00000000";
		ram_buffer(7099) := X"00000000";
		ram_buffer(7100) := X"00000000";
		ram_buffer(7101) := X"00000000";
		ram_buffer(7102) := X"00000000";
		ram_buffer(7103) := X"00000000";
		ram_buffer(7104) := X"00000000";
		ram_buffer(7105) := X"00000000";
		ram_buffer(7106) := X"00000000";
		ram_buffer(7107) := X"00000000";
		ram_buffer(7108) := X"00000000";
		ram_buffer(7109) := X"00000000";
		ram_buffer(7110) := X"00000000";
		ram_buffer(7111) := X"00000000";
		ram_buffer(7112) := X"00000000";
		ram_buffer(7113) := X"00000000";
		ram_buffer(7114) := X"00000000";
		ram_buffer(7115) := X"00000000";
		ram_buffer(7116) := X"00000000";
		ram_buffer(7117) := X"00000000";
		ram_buffer(7118) := X"00000000";
		ram_buffer(7119) := X"00000000";
		ram_buffer(7120) := X"00000000";
		ram_buffer(7121) := X"00000000";
		ram_buffer(7122) := X"00000000";
		ram_buffer(7123) := X"00000000";
		ram_buffer(7124) := X"00000000";
		ram_buffer(7125) := X"00000000";
		ram_buffer(7126) := X"00000000";
		ram_buffer(7127) := X"00000000";
		ram_buffer(7128) := X"00000000";
		ram_buffer(7129) := X"00000000";
		ram_buffer(7130) := X"00000000";
		ram_buffer(7131) := X"00000000";
		ram_buffer(7132) := X"00000000";
		ram_buffer(7133) := X"00000000";
		ram_buffer(7134) := X"00000000";
		ram_buffer(7135) := X"00000000";
		ram_buffer(7136) := X"00000000";
		ram_buffer(7137) := X"00000000";
		ram_buffer(7138) := X"00000000";
		ram_buffer(7139) := X"00000000";
		ram_buffer(7140) := X"00000000";
		ram_buffer(7141) := X"00000000";
		ram_buffer(7142) := X"00000000";
		ram_buffer(7143) := X"00000000";
		ram_buffer(7144) := X"00000000";
		ram_buffer(7145) := X"00000000";
		ram_buffer(7146) := X"00000000";
		ram_buffer(7147) := X"00000000";
		ram_buffer(7148) := X"00000000";
		ram_buffer(7149) := X"00000000";
		ram_buffer(7150) := X"00000000";
		ram_buffer(7151) := X"00000000";
		ram_buffer(7152) := X"00000000";
		ram_buffer(7153) := X"00000000";
		ram_buffer(7154) := X"00000000";
		ram_buffer(7155) := X"00000000";
		ram_buffer(7156) := X"00000000";
		ram_buffer(7157) := X"00000000";
		ram_buffer(7158) := X"00000000";
		ram_buffer(7159) := X"00000000";
		ram_buffer(7160) := X"00000000";
		ram_buffer(7161) := X"00000000";
		ram_buffer(7162) := X"00000000";
		ram_buffer(7163) := X"00000000";
		ram_buffer(7164) := X"00000000";
		ram_buffer(7165) := X"00000000";
		ram_buffer(7166) := X"00000000";
		ram_buffer(7167) := X"00000000";
		ram_buffer(7168) := X"00000000";
		ram_buffer(7169) := X"00000000";
		ram_buffer(7170) := X"00000000";
		ram_buffer(7171) := X"00000000";
		ram_buffer(7172) := X"00000000";
		ram_buffer(7173) := X"00000000";
		ram_buffer(7174) := X"00000000";
		ram_buffer(7175) := X"00000000";
		ram_buffer(7176) := X"00000000";
		ram_buffer(7177) := X"00000000";
		ram_buffer(7178) := X"00000000";
		ram_buffer(7179) := X"00000000";
		ram_buffer(7180) := X"00000000";
		ram_buffer(7181) := X"00000000";
		ram_buffer(7182) := X"00000000";
		ram_buffer(7183) := X"00000000";
		ram_buffer(7184) := X"00000000";
		ram_buffer(7185) := X"00000000";
		ram_buffer(7186) := X"00000000";
		ram_buffer(7187) := X"00000000";
		ram_buffer(7188) := X"00000000";
		ram_buffer(7189) := X"00000000";
		ram_buffer(7190) := X"00000000";
		ram_buffer(7191) := X"00000000";
		ram_buffer(7192) := X"00000000";
		ram_buffer(7193) := X"00000000";
		ram_buffer(7194) := X"00000000";
		ram_buffer(7195) := X"00000000";
		ram_buffer(7196) := X"00000000";
		ram_buffer(7197) := X"00000000";
		ram_buffer(7198) := X"00000000";
		ram_buffer(7199) := X"00000000";
		ram_buffer(7200) := X"00000000";
		ram_buffer(7201) := X"00000000";
		ram_buffer(7202) := X"00000000";
		ram_buffer(7203) := X"00000000";
		ram_buffer(7204) := X"00000000";
		ram_buffer(7205) := X"00000000";
		ram_buffer(7206) := X"00000000";
		ram_buffer(7207) := X"00000000";
		ram_buffer(7208) := X"00000000";
		ram_buffer(7209) := X"00000000";
		ram_buffer(7210) := X"00000000";
		ram_buffer(7211) := X"00000000";
		ram_buffer(7212) := X"00000000";
		ram_buffer(7213) := X"00000000";
		ram_buffer(7214) := X"00000000";
		ram_buffer(7215) := X"00000000";
		ram_buffer(7216) := X"00000000";
		ram_buffer(7217) := X"00000000";
		ram_buffer(7218) := X"00000000";
		ram_buffer(7219) := X"00000000";
		ram_buffer(7220) := X"00000000";
		ram_buffer(7221) := X"00000000";
		ram_buffer(7222) := X"00000000";
		ram_buffer(7223) := X"00000000";
		ram_buffer(7224) := X"00000000";
		ram_buffer(7225) := X"00000000";
		ram_buffer(7226) := X"00000000";
		ram_buffer(7227) := X"00000000";
		ram_buffer(7228) := X"00000000";
		ram_buffer(7229) := X"00000000";
		ram_buffer(7230) := X"00000000";
		ram_buffer(7231) := X"00000000";
		ram_buffer(7232) := X"00000000";
		ram_buffer(7233) := X"00000000";
		ram_buffer(7234) := X"00000000";
		ram_buffer(7235) := X"00000000";
		ram_buffer(7236) := X"00000000";
		ram_buffer(7237) := X"00000000";
		ram_buffer(7238) := X"00000000";
		ram_buffer(7239) := X"00000000";
		ram_buffer(7240) := X"00000000";
		ram_buffer(7241) := X"00000000";
		ram_buffer(7242) := X"00000000";
		ram_buffer(7243) := X"00000000";
		ram_buffer(7244) := X"00000000";
		ram_buffer(7245) := X"00000000";
		ram_buffer(7246) := X"00000000";
		ram_buffer(7247) := X"00000000";
		ram_buffer(7248) := X"00000000";
		ram_buffer(7249) := X"00000000";
		ram_buffer(7250) := X"00000000";
		ram_buffer(7251) := X"00000000";
		ram_buffer(7252) := X"00000000";
		ram_buffer(7253) := X"00000000";
		ram_buffer(7254) := X"00000000";
		ram_buffer(7255) := X"00000000";
		ram_buffer(7256) := X"00000000";
		ram_buffer(7257) := X"00000000";
		ram_buffer(7258) := X"00000000";
		ram_buffer(7259) := X"00000000";
		ram_buffer(7260) := X"00000000";
		ram_buffer(7261) := X"00000000";
		ram_buffer(7262) := X"00000000";
		ram_buffer(7263) := X"00000000";
		ram_buffer(7264) := X"00000000";
		ram_buffer(7265) := X"00000000";
		ram_buffer(7266) := X"00000000";
		ram_buffer(7267) := X"00000000";
		ram_buffer(7268) := X"00000000";
		ram_buffer(7269) := X"00000000";
		ram_buffer(7270) := X"00000000";
		ram_buffer(7271) := X"00000000";
		ram_buffer(7272) := X"00000000";
		ram_buffer(7273) := X"00000000";
		ram_buffer(7274) := X"00000000";
		ram_buffer(7275) := X"00000000";
		ram_buffer(7276) := X"00000000";
		ram_buffer(7277) := X"00000000";
		ram_buffer(7278) := X"00000000";
		ram_buffer(7279) := X"00000000";
		ram_buffer(7280) := X"00000000";
		ram_buffer(7281) := X"00000000";
		ram_buffer(7282) := X"00000000";
		ram_buffer(7283) := X"00000000";
		ram_buffer(7284) := X"00000000";
		ram_buffer(7285) := X"00000000";
		ram_buffer(7286) := X"00000000";
		ram_buffer(7287) := X"00000000";
		ram_buffer(7288) := X"00000000";
		ram_buffer(7289) := X"00000000";
		ram_buffer(7290) := X"00000000";
		ram_buffer(7291) := X"00000000";
		ram_buffer(7292) := X"00000000";
		ram_buffer(7293) := X"00000000";
		ram_buffer(7294) := X"00000000";
		ram_buffer(7295) := X"00000000";
		ram_buffer(7296) := X"00000000";
		ram_buffer(7297) := X"00000000";
		ram_buffer(7298) := X"00000000";
		ram_buffer(7299) := X"00000000";
		ram_buffer(7300) := X"00000000";
		ram_buffer(7301) := X"00000000";
		ram_buffer(7302) := X"00000000";
		ram_buffer(7303) := X"00000000";
		ram_buffer(7304) := X"00000000";
		ram_buffer(7305) := X"00000000";
		ram_buffer(7306) := X"00000000";
		ram_buffer(7307) := X"00000000";
		ram_buffer(7308) := X"00000000";
		ram_buffer(7309) := X"00000000";
		ram_buffer(7310) := X"00000000";
		ram_buffer(7311) := X"00000000";
		ram_buffer(7312) := X"00000000";
		ram_buffer(7313) := X"00000000";
		ram_buffer(7314) := X"00000000";
		ram_buffer(7315) := X"00000000";
		ram_buffer(7316) := X"00000000";
		ram_buffer(7317) := X"00000000";
		ram_buffer(7318) := X"00000000";
		ram_buffer(7319) := X"00000000";
		ram_buffer(7320) := X"00000000";
		ram_buffer(7321) := X"00000000";
		ram_buffer(7322) := X"00000000";
		ram_buffer(7323) := X"00000000";
		ram_buffer(7324) := X"00000000";
		ram_buffer(7325) := X"00000000";
		ram_buffer(7326) := X"00000000";
		ram_buffer(7327) := X"00000000";
		ram_buffer(7328) := X"00000000";
		ram_buffer(7329) := X"00000000";
		ram_buffer(7330) := X"00000000";
		ram_buffer(7331) := X"00000000";
		ram_buffer(7332) := X"00000000";
		ram_buffer(7333) := X"00000000";
		ram_buffer(7334) := X"00000000";
		ram_buffer(7335) := X"00000000";
		ram_buffer(7336) := X"00000000";
		ram_buffer(7337) := X"00000000";
		ram_buffer(7338) := X"00000000";
		ram_buffer(7339) := X"00000000";
		ram_buffer(7340) := X"00000000";
		ram_buffer(7341) := X"00000000";
		ram_buffer(7342) := X"00000000";
		ram_buffer(7343) := X"00000000";
		ram_buffer(7344) := X"00000000";
		ram_buffer(7345) := X"00000000";
		ram_buffer(7346) := X"00000000";
		ram_buffer(7347) := X"00000000";
		ram_buffer(7348) := X"00000000";
		ram_buffer(7349) := X"00000000";
		ram_buffer(7350) := X"00000000";
		ram_buffer(7351) := X"00000000";
		ram_buffer(7352) := X"00000000";
		ram_buffer(7353) := X"00000000";
		ram_buffer(7354) := X"00000000";
		ram_buffer(7355) := X"00000000";
		ram_buffer(7356) := X"00000000";
		ram_buffer(7357) := X"00000000";
		ram_buffer(7358) := X"00000000";
		ram_buffer(7359) := X"00000000";
		ram_buffer(7360) := X"00000000";
		ram_buffer(7361) := X"00000000";
		ram_buffer(7362) := X"00000000";
		ram_buffer(7363) := X"00000000";
		ram_buffer(7364) := X"00000000";
		ram_buffer(7365) := X"00000000";
		ram_buffer(7366) := X"00000000";
		ram_buffer(7367) := X"00000000";
		ram_buffer(7368) := X"00000000";
		ram_buffer(7369) := X"00000000";
		ram_buffer(7370) := X"00000000";
		ram_buffer(7371) := X"00000000";
		ram_buffer(7372) := X"00000000";
		ram_buffer(7373) := X"00000000";
		ram_buffer(7374) := X"00000000";
		ram_buffer(7375) := X"00000000";
		ram_buffer(7376) := X"00000000";
		ram_buffer(7377) := X"00000000";
		ram_buffer(7378) := X"00000000";
		ram_buffer(7379) := X"00000000";
		ram_buffer(7380) := X"00000000";
		ram_buffer(7381) := X"00000000";
		ram_buffer(7382) := X"00000000";
		ram_buffer(7383) := X"00000000";
		ram_buffer(7384) := X"00000000";
		ram_buffer(7385) := X"00000000";
		ram_buffer(7386) := X"00000000";
		ram_buffer(7387) := X"00000000";
		ram_buffer(7388) := X"00000000";
		ram_buffer(7389) := X"00000000";
		ram_buffer(7390) := X"00000000";
		ram_buffer(7391) := X"00000000";
		ram_buffer(7392) := X"00000000";
		ram_buffer(7393) := X"00000000";
		ram_buffer(7394) := X"00000000";
		ram_buffer(7395) := X"00000000";
		ram_buffer(7396) := X"00000000";
		ram_buffer(7397) := X"00000000";
		ram_buffer(7398) := X"00000000";
		ram_buffer(7399) := X"00000000";
		ram_buffer(7400) := X"00000000";
		ram_buffer(7401) := X"00000000";
		ram_buffer(7402) := X"00000000";
		ram_buffer(7403) := X"00000000";
		ram_buffer(7404) := X"00000000";
		ram_buffer(7405) := X"00000000";
		ram_buffer(7406) := X"00000000";
		ram_buffer(7407) := X"00000000";
		ram_buffer(7408) := X"00000000";
		ram_buffer(7409) := X"00000000";
		ram_buffer(7410) := X"00000000";
		ram_buffer(7411) := X"00000000";
		ram_buffer(7412) := X"00000000";
		ram_buffer(7413) := X"00000000";
		ram_buffer(7414) := X"00000000";
		ram_buffer(7415) := X"00000000";
		ram_buffer(7416) := X"00000000";
		ram_buffer(7417) := X"00000000";
		ram_buffer(7418) := X"00000000";
		ram_buffer(7419) := X"00000000";
		ram_buffer(7420) := X"00000000";
		ram_buffer(7421) := X"00000000";
		ram_buffer(7422) := X"00000000";
		ram_buffer(7423) := X"00000000";
		ram_buffer(7424) := X"00000000";
		ram_buffer(7425) := X"00000000";
		ram_buffer(7426) := X"00000000";
		ram_buffer(7427) := X"00000000";
		ram_buffer(7428) := X"00000000";
		ram_buffer(7429) := X"00000000";
		ram_buffer(7430) := X"00000000";
		ram_buffer(7431) := X"00000000";
		ram_buffer(7432) := X"00000000";
		ram_buffer(7433) := X"00000000";
		ram_buffer(7434) := X"00000000";
		ram_buffer(7435) := X"00000000";
		ram_buffer(7436) := X"00000000";
		ram_buffer(7437) := X"00000000";
		ram_buffer(7438) := X"00000000";
		ram_buffer(7439) := X"00000000";
		ram_buffer(7440) := X"00000000";
		ram_buffer(7441) := X"00000000";
		ram_buffer(7442) := X"00000000";
		ram_buffer(7443) := X"00000000";
		ram_buffer(7444) := X"00000000";
		ram_buffer(7445) := X"00000000";
		ram_buffer(7446) := X"00000000";
		ram_buffer(7447) := X"00000000";
		ram_buffer(7448) := X"00000000";
		ram_buffer(7449) := X"00000000";
		ram_buffer(7450) := X"00000000";
		ram_buffer(7451) := X"00000000";
		ram_buffer(7452) := X"00000000";
		ram_buffer(7453) := X"00000000";
		ram_buffer(7454) := X"00000000";
		ram_buffer(7455) := X"00000000";
		ram_buffer(7456) := X"00000000";
		ram_buffer(7457) := X"00000000";
		ram_buffer(7458) := X"00000000";
		ram_buffer(7459) := X"00000000";
		ram_buffer(7460) := X"00000000";
		ram_buffer(7461) := X"00000000";
		ram_buffer(7462) := X"00000000";
		ram_buffer(7463) := X"00000000";
		ram_buffer(7464) := X"00000000";
		ram_buffer(7465) := X"00000000";
		ram_buffer(7466) := X"00000000";
		ram_buffer(7467) := X"00000000";
		ram_buffer(7468) := X"00000000";
		ram_buffer(7469) := X"00000000";
		ram_buffer(7470) := X"00000000";
		ram_buffer(7471) := X"00000000";
		ram_buffer(7472) := X"00000000";
		ram_buffer(7473) := X"00000000";
		ram_buffer(7474) := X"00000000";
		ram_buffer(7475) := X"00000000";
		ram_buffer(7476) := X"00000000";
		ram_buffer(7477) := X"00000000";
		ram_buffer(7478) := X"00000000";
		ram_buffer(7479) := X"00000000";
		ram_buffer(7480) := X"00000000";
		ram_buffer(7481) := X"00000000";
		ram_buffer(7482) := X"00000000";
		ram_buffer(7483) := X"00000000";
		ram_buffer(7484) := X"00000000";
		ram_buffer(7485) := X"00000000";
		ram_buffer(7486) := X"00000000";
		ram_buffer(7487) := X"00000000";
		ram_buffer(7488) := X"00000000";
		ram_buffer(7489) := X"00000000";
		ram_buffer(7490) := X"00000000";
		ram_buffer(7491) := X"00000000";
		ram_buffer(7492) := X"00000000";
		ram_buffer(7493) := X"00000000";
		ram_buffer(7494) := X"00000000";
		ram_buffer(7495) := X"00000000";
		ram_buffer(7496) := X"00000000";
		ram_buffer(7497) := X"00000000";
		ram_buffer(7498) := X"00000000";
		ram_buffer(7499) := X"00000000";
		ram_buffer(7500) := X"00000000";
		ram_buffer(7501) := X"00000000";
		ram_buffer(7502) := X"00000000";
		ram_buffer(7503) := X"00000000";
		ram_buffer(7504) := X"00000000";
		ram_buffer(7505) := X"00000000";
		ram_buffer(7506) := X"00000000";
		ram_buffer(7507) := X"00000000";
		ram_buffer(7508) := X"00000000";
		ram_buffer(7509) := X"00000000";
		ram_buffer(7510) := X"00000000";
		ram_buffer(7511) := X"00000000";
		ram_buffer(7512) := X"00000000";
		ram_buffer(7513) := X"00000000";
		ram_buffer(7514) := X"00000000";
		ram_buffer(7515) := X"00000000";
		ram_buffer(7516) := X"00000000";
		ram_buffer(7517) := X"00000000";
		ram_buffer(7518) := X"00000000";
		ram_buffer(7519) := X"00000000";
		ram_buffer(7520) := X"00000000";
		ram_buffer(7521) := X"00000000";
		ram_buffer(7522) := X"00000000";
		ram_buffer(7523) := X"00000000";
		ram_buffer(7524) := X"00000000";
		ram_buffer(7525) := X"00000000";
		ram_buffer(7526) := X"00000000";
		ram_buffer(7527) := X"00000000";
		ram_buffer(7528) := X"00000000";
		ram_buffer(7529) := X"00000000";
		ram_buffer(7530) := X"00000000";
		ram_buffer(7531) := X"00000000";
		ram_buffer(7532) := X"00000000";
		ram_buffer(7533) := X"00000000";
		ram_buffer(7534) := X"00000000";
		ram_buffer(7535) := X"00000000";
		ram_buffer(7536) := X"00000000";
		ram_buffer(7537) := X"00000000";
		ram_buffer(7538) := X"00000000";
		ram_buffer(7539) := X"00000000";
		ram_buffer(7540) := X"00000000";
		ram_buffer(7541) := X"00000000";
		ram_buffer(7542) := X"00000000";
		ram_buffer(7543) := X"00000000";
		ram_buffer(7544) := X"00000000";
		ram_buffer(7545) := X"00000000";
		ram_buffer(7546) := X"00000000";
		ram_buffer(7547) := X"00000000";
		ram_buffer(7548) := X"00000000";
		ram_buffer(7549) := X"00000000";
		ram_buffer(7550) := X"00000000";
		ram_buffer(7551) := X"00000000";
		ram_buffer(7552) := X"00000000";
		ram_buffer(7553) := X"00000000";
		ram_buffer(7554) := X"00000000";
		ram_buffer(7555) := X"00000000";
		ram_buffer(7556) := X"00000000";
		ram_buffer(7557) := X"00000000";
		ram_buffer(7558) := X"00000000";
		ram_buffer(7559) := X"00000000";
		ram_buffer(7560) := X"00000000";
		ram_buffer(7561) := X"00000000";
		ram_buffer(7562) := X"00000000";
		ram_buffer(7563) := X"00000000";
		ram_buffer(7564) := X"00000000";
		ram_buffer(7565) := X"00000000";
		ram_buffer(7566) := X"00000000";
		ram_buffer(7567) := X"00000000";
		ram_buffer(7568) := X"00000000";
		ram_buffer(7569) := X"00000000";
		ram_buffer(7570) := X"00000000";
		ram_buffer(7571) := X"00000000";
		ram_buffer(7572) := X"00000000";
		ram_buffer(7573) := X"00000000";
		ram_buffer(7574) := X"00000000";
		ram_buffer(7575) := X"00000000";
		ram_buffer(7576) := X"00000000";
		ram_buffer(7577) := X"00000000";
		ram_buffer(7578) := X"00000000";
		ram_buffer(7579) := X"00000000";
		ram_buffer(7580) := X"00000000";
		ram_buffer(7581) := X"00000000";
		ram_buffer(7582) := X"00000000";
		ram_buffer(7583) := X"00000000";
		ram_buffer(7584) := X"00000000";
		ram_buffer(7585) := X"00000000";
		ram_buffer(7586) := X"00000000";
		ram_buffer(7587) := X"00000000";
		ram_buffer(7588) := X"00000000";
		ram_buffer(7589) := X"00000000";
		ram_buffer(7590) := X"00000000";
		ram_buffer(7591) := X"00000000";
		ram_buffer(7592) := X"00000000";
		ram_buffer(7593) := X"00000000";
		ram_buffer(7594) := X"00000000";
		ram_buffer(7595) := X"00000000";
		ram_buffer(7596) := X"00000000";
		ram_buffer(7597) := X"00000000";
		ram_buffer(7598) := X"00000000";
		ram_buffer(7599) := X"00000000";
		ram_buffer(7600) := X"00000000";
		ram_buffer(7601) := X"00000000";
		ram_buffer(7602) := X"00000000";
		ram_buffer(7603) := X"00000000";
		ram_buffer(7604) := X"00000000";
		ram_buffer(7605) := X"00000000";
		ram_buffer(7606) := X"00000000";
		ram_buffer(7607) := X"00000000";
		ram_buffer(7608) := X"00000000";
		ram_buffer(7609) := X"00000000";
		ram_buffer(7610) := X"00000000";
		ram_buffer(7611) := X"00000000";
		ram_buffer(7612) := X"00000000";
		ram_buffer(7613) := X"00000000";
		ram_buffer(7614) := X"00000000";
		ram_buffer(7615) := X"00000000";
		ram_buffer(7616) := X"00000000";
		ram_buffer(7617) := X"00000000";
		ram_buffer(7618) := X"00000000";
		ram_buffer(7619) := X"00000000";
		ram_buffer(7620) := X"00000000";
		ram_buffer(7621) := X"00000000";
		ram_buffer(7622) := X"00000000";
		ram_buffer(7623) := X"00000000";
		ram_buffer(7624) := X"00000000";
		ram_buffer(7625) := X"00000000";
		ram_buffer(7626) := X"00000000";
		ram_buffer(7627) := X"00000000";
		ram_buffer(7628) := X"00000000";
		ram_buffer(7629) := X"00000000";
		ram_buffer(7630) := X"00000000";
		ram_buffer(7631) := X"00000000";
		ram_buffer(7632) := X"00000000";
		ram_buffer(7633) := X"00000000";
		ram_buffer(7634) := X"00000000";
		ram_buffer(7635) := X"00000000";
		ram_buffer(7636) := X"00000000";
		ram_buffer(7637) := X"00000000";
		ram_buffer(7638) := X"00000000";
		ram_buffer(7639) := X"00000000";
		ram_buffer(7640) := X"00000000";
		ram_buffer(7641) := X"00000000";
		ram_buffer(7642) := X"00000000";
		ram_buffer(7643) := X"00000000";
		ram_buffer(7644) := X"00000000";
		ram_buffer(7645) := X"00000000";
		ram_buffer(7646) := X"00000000";
		ram_buffer(7647) := X"00000000";
		ram_buffer(7648) := X"00000000";
		ram_buffer(7649) := X"00000000";
		ram_buffer(7650) := X"00000000";
		ram_buffer(7651) := X"00000000";
		ram_buffer(7652) := X"00000000";
		ram_buffer(7653) := X"00000000";
		ram_buffer(7654) := X"00000000";
		ram_buffer(7655) := X"00000000";
		ram_buffer(7656) := X"00000000";
		ram_buffer(7657) := X"00000000";
		ram_buffer(7658) := X"00000000";
		ram_buffer(7659) := X"00000000";
		ram_buffer(7660) := X"00000000";
		ram_buffer(7661) := X"00000000";
		ram_buffer(7662) := X"00000000";
		ram_buffer(7663) := X"00000000";
		ram_buffer(7664) := X"00000000";
		ram_buffer(7665) := X"00000000";
		ram_buffer(7666) := X"00000000";
		ram_buffer(7667) := X"00000000";
		ram_buffer(7668) := X"00000000";
		ram_buffer(7669) := X"00000000";
		ram_buffer(7670) := X"00000000";
		ram_buffer(7671) := X"00000000";
		ram_buffer(7672) := X"00000000";
		ram_buffer(7673) := X"00000000";
		ram_buffer(7674) := X"00000000";
		ram_buffer(7675) := X"00000000";
		ram_buffer(7676) := X"00000000";
		ram_buffer(7677) := X"00000000";
		ram_buffer(7678) := X"00000000";
		ram_buffer(7679) := X"00000000";
		ram_buffer(7680) := X"00000000";
		ram_buffer(7681) := X"00000000";
		ram_buffer(7682) := X"00000000";
		ram_buffer(7683) := X"00000000";
		ram_buffer(7684) := X"00000000";
		ram_buffer(7685) := X"00000000";
		ram_buffer(7686) := X"00000000";
		ram_buffer(7687) := X"00000000";
		ram_buffer(7688) := X"00000000";
		ram_buffer(7689) := X"00000000";
		ram_buffer(7690) := X"00000000";
		ram_buffer(7691) := X"00000000";
		ram_buffer(7692) := X"00000000";
		ram_buffer(7693) := X"00000000";
		ram_buffer(7694) := X"00000000";
		ram_buffer(7695) := X"00000000";
		ram_buffer(7696) := X"00000000";
		ram_buffer(7697) := X"00000000";
		ram_buffer(7698) := X"00000000";
		ram_buffer(7699) := X"00000000";
		ram_buffer(7700) := X"00000000";
		ram_buffer(7701) := X"00000000";
		ram_buffer(7702) := X"00000000";
		ram_buffer(7703) := X"00000000";
		ram_buffer(7704) := X"00000000";
		ram_buffer(7705) := X"00000000";
		ram_buffer(7706) := X"00000000";
		ram_buffer(7707) := X"00000000";
		ram_buffer(7708) := X"00000000";
		ram_buffer(7709) := X"00000000";
		ram_buffer(7710) := X"00000000";
		ram_buffer(7711) := X"00000000";
		ram_buffer(7712) := X"00000000";
		ram_buffer(7713) := X"00000000";
		ram_buffer(7714) := X"00000000";
		ram_buffer(7715) := X"00000000";
		ram_buffer(7716) := X"00000000";
		ram_buffer(7717) := X"00000000";
		ram_buffer(7718) := X"00000000";
		ram_buffer(7719) := X"00000000";
		ram_buffer(7720) := X"00000000";
		ram_buffer(7721) := X"00000000";
		ram_buffer(7722) := X"00000000";
		ram_buffer(7723) := X"00000000";
		ram_buffer(7724) := X"00000000";
		ram_buffer(7725) := X"00000000";
		ram_buffer(7726) := X"00000000";
		ram_buffer(7727) := X"00000000";
		ram_buffer(7728) := X"00000000";
		ram_buffer(7729) := X"00000000";
		ram_buffer(7730) := X"00000000";
		ram_buffer(7731) := X"00000000";
		ram_buffer(7732) := X"00000000";
		ram_buffer(7733) := X"00000000";
		ram_buffer(7734) := X"00000000";
		ram_buffer(7735) := X"00000000";
		ram_buffer(7736) := X"00000000";
		ram_buffer(7737) := X"00000000";
		ram_buffer(7738) := X"00000000";
		ram_buffer(7739) := X"00000000";
		ram_buffer(7740) := X"00000000";
		ram_buffer(7741) := X"00000000";
		ram_buffer(7742) := X"00000000";
		ram_buffer(7743) := X"00000000";
		ram_buffer(7744) := X"00000000";
		ram_buffer(7745) := X"00000000";
		ram_buffer(7746) := X"00000000";
		ram_buffer(7747) := X"00000000";
		ram_buffer(7748) := X"00000000";
		ram_buffer(7749) := X"00000000";
		ram_buffer(7750) := X"00000000";
		ram_buffer(7751) := X"00000000";
		ram_buffer(7752) := X"00000000";
		ram_buffer(7753) := X"00000000";
		ram_buffer(7754) := X"00000000";
		ram_buffer(7755) := X"00000000";
		ram_buffer(7756) := X"00000000";
		ram_buffer(7757) := X"00000000";
		ram_buffer(7758) := X"00000000";
		ram_buffer(7759) := X"00000000";
		ram_buffer(7760) := X"00000000";
		ram_buffer(7761) := X"00000000";
		ram_buffer(7762) := X"00000000";
		ram_buffer(7763) := X"00000000";
		ram_buffer(7764) := X"00000000";
		ram_buffer(7765) := X"00000000";
		ram_buffer(7766) := X"00000000";
		ram_buffer(7767) := X"00000000";
		ram_buffer(7768) := X"00000000";
		ram_buffer(7769) := X"00000000";
		ram_buffer(7770) := X"00000000";
		ram_buffer(7771) := X"00000000";
		ram_buffer(7772) := X"00000000";
		ram_buffer(7773) := X"00000000";
		ram_buffer(7774) := X"00000000";
		ram_buffer(7775) := X"00000000";
		ram_buffer(7776) := X"00000000";
		ram_buffer(7777) := X"00000000";
		ram_buffer(7778) := X"00000000";
		ram_buffer(7779) := X"00000000";
		ram_buffer(7780) := X"00000000";
		ram_buffer(7781) := X"00000000";
		ram_buffer(7782) := X"00000000";
		ram_buffer(7783) := X"00000000";
		ram_buffer(7784) := X"00000000";
		ram_buffer(7785) := X"00000000";
		ram_buffer(7786) := X"00000000";
		ram_buffer(7787) := X"00000000";
		ram_buffer(7788) := X"00000000";
		ram_buffer(7789) := X"00000000";
		ram_buffer(7790) := X"00000000";
		ram_buffer(7791) := X"00000000";
		ram_buffer(7792) := X"00000000";
		ram_buffer(7793) := X"00000000";
		ram_buffer(7794) := X"00000000";
		ram_buffer(7795) := X"00000000";
		ram_buffer(7796) := X"00000000";
		ram_buffer(7797) := X"00000000";
		ram_buffer(7798) := X"00000000";
		ram_buffer(7799) := X"00000000";
		ram_buffer(7800) := X"00000000";
		ram_buffer(7801) := X"00000000";
		ram_buffer(7802) := X"00000000";
		ram_buffer(7803) := X"00000000";
		ram_buffer(7804) := X"00000000";
		ram_buffer(7805) := X"00000000";
		ram_buffer(7806) := X"00000000";
		ram_buffer(7807) := X"00000000";
		ram_buffer(7808) := X"00000000";
		ram_buffer(7809) := X"00000000";
		ram_buffer(7810) := X"00000000";
		ram_buffer(7811) := X"00000000";
		ram_buffer(7812) := X"00000000";
		ram_buffer(7813) := X"00000000";
		ram_buffer(7814) := X"00000000";
		ram_buffer(7815) := X"00000000";
		ram_buffer(7816) := X"00000000";
		ram_buffer(7817) := X"00000000";
		ram_buffer(7818) := X"00000000";
		ram_buffer(7819) := X"00000000";
		ram_buffer(7820) := X"00000000";
		ram_buffer(7821) := X"00000000";
		ram_buffer(7822) := X"00000000";
		ram_buffer(7823) := X"00000000";
		ram_buffer(7824) := X"00000000";
		ram_buffer(7825) := X"00000000";
		ram_buffer(7826) := X"00000000";
		ram_buffer(7827) := X"00000000";
		ram_buffer(7828) := X"00000000";
		ram_buffer(7829) := X"00000000";
		ram_buffer(7830) := X"00000000";
		ram_buffer(7831) := X"00000000";
		ram_buffer(7832) := X"00000000";
		ram_buffer(7833) := X"00000000";
		ram_buffer(7834) := X"00000000";
		ram_buffer(7835) := X"00000000";
		ram_buffer(7836) := X"00000000";
		ram_buffer(7837) := X"00000000";
		ram_buffer(7838) := X"00000000";
		ram_buffer(7839) := X"00000000";
		ram_buffer(7840) := X"00000000";
		ram_buffer(7841) := X"00000000";
		ram_buffer(7842) := X"00000000";
		ram_buffer(7843) := X"00000000";
		ram_buffer(7844) := X"00000000";
		ram_buffer(7845) := X"00000000";
		ram_buffer(7846) := X"00000000";
		ram_buffer(7847) := X"00000000";
		ram_buffer(7848) := X"00000000";
		ram_buffer(7849) := X"00000000";
		ram_buffer(7850) := X"00000000";
		ram_buffer(7851) := X"00000000";
		ram_buffer(7852) := X"00000000";
		ram_buffer(7853) := X"00000000";
		ram_buffer(7854) := X"00000000";
		ram_buffer(7855) := X"00000000";
		ram_buffer(7856) := X"00000000";
		ram_buffer(7857) := X"00000000";
		ram_buffer(7858) := X"00000000";
		ram_buffer(7859) := X"00000000";
		ram_buffer(7860) := X"00000000";
		ram_buffer(7861) := X"00000000";
		ram_buffer(7862) := X"00000000";
		ram_buffer(7863) := X"00000000";
		ram_buffer(7864) := X"00000000";
		ram_buffer(7865) := X"00000000";
		ram_buffer(7866) := X"00000000";
		ram_buffer(7867) := X"00000000";
		ram_buffer(7868) := X"00000000";
		ram_buffer(7869) := X"00000000";
		ram_buffer(7870) := X"00000000";
		ram_buffer(7871) := X"00000000";
		ram_buffer(7872) := X"00000000";
		ram_buffer(7873) := X"00000000";
		ram_buffer(7874) := X"00000000";
		ram_buffer(7875) := X"00000000";
		ram_buffer(7876) := X"00000000";
		ram_buffer(7877) := X"00000000";
		ram_buffer(7878) := X"00000000";
		ram_buffer(7879) := X"00000000";
		ram_buffer(7880) := X"00000000";
		ram_buffer(7881) := X"00000000";
		ram_buffer(7882) := X"00000000";
		ram_buffer(7883) := X"00000000";
		ram_buffer(7884) := X"00000000";
		ram_buffer(7885) := X"00000000";
		ram_buffer(7886) := X"00000000";
		ram_buffer(7887) := X"00000000";
		ram_buffer(7888) := X"00000000";
		ram_buffer(7889) := X"00000000";
		ram_buffer(7890) := X"00000000";
		ram_buffer(7891) := X"00000000";
		ram_buffer(7892) := X"00000000";
		ram_buffer(7893) := X"00000000";
		ram_buffer(7894) := X"00000000";
		ram_buffer(7895) := X"00000000";
		ram_buffer(7896) := X"00000000";
		ram_buffer(7897) := X"00000000";
		ram_buffer(7898) := X"00000000";
		ram_buffer(7899) := X"00000000";
		ram_buffer(7900) := X"00000000";
		ram_buffer(7901) := X"00000000";
		ram_buffer(7902) := X"00000000";
		ram_buffer(7903) := X"00000000";
		ram_buffer(7904) := X"00000000";
		ram_buffer(7905) := X"00000000";
		ram_buffer(7906) := X"00000000";
		ram_buffer(7907) := X"00000000";
		ram_buffer(7908) := X"00000000";
		ram_buffer(7909) := X"00000000";
		ram_buffer(7910) := X"00000000";
		ram_buffer(7911) := X"00000000";
		ram_buffer(7912) := X"00000000";
		ram_buffer(7913) := X"00000000";
		ram_buffer(7914) := X"00000000";
		ram_buffer(7915) := X"00000000";
		ram_buffer(7916) := X"00000000";
		ram_buffer(7917) := X"00000000";
		ram_buffer(7918) := X"00000000";
		ram_buffer(7919) := X"00000000";
		ram_buffer(7920) := X"00000000";
		ram_buffer(7921) := X"00000000";
		ram_buffer(7922) := X"00000000";
		ram_buffer(7923) := X"00000000";
		ram_buffer(7924) := X"00000000";
		ram_buffer(7925) := X"00000000";
		ram_buffer(7926) := X"00000000";
		ram_buffer(7927) := X"00000000";
		ram_buffer(7928) := X"00000000";
		ram_buffer(7929) := X"00000000";
		ram_buffer(7930) := X"00000000";
		ram_buffer(7931) := X"00000000";
		ram_buffer(7932) := X"00000000";
		ram_buffer(7933) := X"00000000";
		ram_buffer(7934) := X"00000000";
		ram_buffer(7935) := X"00000000";
		ram_buffer(7936) := X"00000000";
		ram_buffer(7937) := X"00000000";
		ram_buffer(7938) := X"00000000";
		ram_buffer(7939) := X"00000000";
		ram_buffer(7940) := X"00000000";
		ram_buffer(7941) := X"00000000";
		ram_buffer(7942) := X"00000000";
		ram_buffer(7943) := X"00000000";
		ram_buffer(7944) := X"00000000";
		ram_buffer(7945) := X"00000000";
		ram_buffer(7946) := X"00000000";
		ram_buffer(7947) := X"00000000";
		ram_buffer(7948) := X"00000000";
		ram_buffer(7949) := X"00000000";
		ram_buffer(7950) := X"00000000";
		ram_buffer(7951) := X"00000000";
		ram_buffer(7952) := X"00000000";
		ram_buffer(7953) := X"00000000";
		ram_buffer(7954) := X"00000000";
		ram_buffer(7955) := X"00000000";
		ram_buffer(7956) := X"00000000";
		ram_buffer(7957) := X"00000000";
		ram_buffer(7958) := X"00000000";
		ram_buffer(7959) := X"00000000";
		ram_buffer(7960) := X"00000000";
		ram_buffer(7961) := X"00000000";
		ram_buffer(7962) := X"00000000";
		ram_buffer(7963) := X"00000000";
		ram_buffer(7964) := X"00000000";
		ram_buffer(7965) := X"00000000";
		ram_buffer(7966) := X"00000000";
		ram_buffer(7967) := X"00000000";
		ram_buffer(7968) := X"00000000";
		ram_buffer(7969) := X"00000000";
		ram_buffer(7970) := X"00000000";
		ram_buffer(7971) := X"00000000";
		ram_buffer(7972) := X"00000000";
		ram_buffer(7973) := X"00000000";
		ram_buffer(7974) := X"00000000";
		ram_buffer(7975) := X"00000000";
		ram_buffer(7976) := X"00000000";
		ram_buffer(7977) := X"00000000";
		ram_buffer(7978) := X"00000000";
		ram_buffer(7979) := X"00000000";
		ram_buffer(7980) := X"00000000";
		ram_buffer(7981) := X"00000000";
		ram_buffer(7982) := X"00000000";
		ram_buffer(7983) := X"00000000";
		ram_buffer(7984) := X"00000000";
		ram_buffer(7985) := X"00000000";
		ram_buffer(7986) := X"00000000";
		ram_buffer(7987) := X"00000000";
		ram_buffer(7988) := X"00000000";
		ram_buffer(7989) := X"00000000";
		ram_buffer(7990) := X"00000000";
		ram_buffer(7991) := X"00000000";
		ram_buffer(7992) := X"00000000";
		ram_buffer(7993) := X"00000000";
		ram_buffer(7994) := X"00000000";
		ram_buffer(7995) := X"00000000";
		ram_buffer(7996) := X"00000000";
		ram_buffer(7997) := X"00000000";
		ram_buffer(7998) := X"00000000";
		ram_buffer(7999) := X"00000000";
		ram_buffer(8000) := X"00000000";
		ram_buffer(8001) := X"00000000";
		ram_buffer(8002) := X"00000000";
		ram_buffer(8003) := X"00000000";
		ram_buffer(8004) := X"00000000";
		ram_buffer(8005) := X"00000000";
		ram_buffer(8006) := X"00000000";
		ram_buffer(8007) := X"00000000";
		ram_buffer(8008) := X"00000000";
		ram_buffer(8009) := X"00000000";
		ram_buffer(8010) := X"00000000";
		ram_buffer(8011) := X"00000000";
		ram_buffer(8012) := X"00000000";
		ram_buffer(8013) := X"00000000";
		ram_buffer(8014) := X"00000000";
		ram_buffer(8015) := X"00000000";
		ram_buffer(8016) := X"00000000";
		ram_buffer(8017) := X"00000000";
		ram_buffer(8018) := X"00000000";
		ram_buffer(8019) := X"00000000";
		ram_buffer(8020) := X"00000000";
		ram_buffer(8021) := X"00000000";
		ram_buffer(8022) := X"00000000";
		ram_buffer(8023) := X"00000000";
		ram_buffer(8024) := X"00000000";
		ram_buffer(8025) := X"00000000";
		ram_buffer(8026) := X"00000000";
		ram_buffer(8027) := X"00000000";
		ram_buffer(8028) := X"00000000";
		ram_buffer(8029) := X"00000000";
		ram_buffer(8030) := X"00000000";
		ram_buffer(8031) := X"00000000";
		ram_buffer(8032) := X"00000000";
		ram_buffer(8033) := X"00000000";
		ram_buffer(8034) := X"00000000";
		ram_buffer(8035) := X"00000000";
		ram_buffer(8036) := X"00000000";
		ram_buffer(8037) := X"00000000";
		ram_buffer(8038) := X"00000000";
		ram_buffer(8039) := X"00000000";
		ram_buffer(8040) := X"00000000";
		ram_buffer(8041) := X"00000000";
		ram_buffer(8042) := X"00000000";
		ram_buffer(8043) := X"00000000";
		ram_buffer(8044) := X"00000000";
		ram_buffer(8045) := X"00000000";
		ram_buffer(8046) := X"00000000";
		ram_buffer(8047) := X"00000000";
		ram_buffer(8048) := X"00000000";
		ram_buffer(8049) := X"00000000";
		ram_buffer(8050) := X"00000000";
		ram_buffer(8051) := X"00000000";
		ram_buffer(8052) := X"00000000";
		ram_buffer(8053) := X"00000000";
		ram_buffer(8054) := X"00000000";
		ram_buffer(8055) := X"00000000";
		ram_buffer(8056) := X"00000000";
		ram_buffer(8057) := X"00000000";
		ram_buffer(8058) := X"00000000";
		ram_buffer(8059) := X"00000000";
		ram_buffer(8060) := X"00000000";
		ram_buffer(8061) := X"00000000";
		ram_buffer(8062) := X"00000000";
		ram_buffer(8063) := X"00000000";
		ram_buffer(8064) := X"00000000";
		ram_buffer(8065) := X"00000000";
		ram_buffer(8066) := X"00000000";
		ram_buffer(8067) := X"00000000";
		ram_buffer(8068) := X"00000000";
		ram_buffer(8069) := X"00000000";
		ram_buffer(8070) := X"00000000";
		ram_buffer(8071) := X"00000000";
		ram_buffer(8072) := X"00000000";
		ram_buffer(8073) := X"00000000";
		ram_buffer(8074) := X"00000000";
		ram_buffer(8075) := X"00000000";
		ram_buffer(8076) := X"00000000";
		ram_buffer(8077) := X"00000000";
		ram_buffer(8078) := X"00000000";
		ram_buffer(8079) := X"00000000";
		ram_buffer(8080) := X"00000000";
		ram_buffer(8081) := X"00000000";
		ram_buffer(8082) := X"00000000";
		ram_buffer(8083) := X"00000000";
		ram_buffer(8084) := X"00000000";
		ram_buffer(8085) := X"00000000";
		ram_buffer(8086) := X"00000000";
		ram_buffer(8087) := X"00000000";
		ram_buffer(8088) := X"00000000";
		ram_buffer(8089) := X"00000000";
		ram_buffer(8090) := X"00000000";
		ram_buffer(8091) := X"00000000";
		ram_buffer(8092) := X"00000000";
		ram_buffer(8093) := X"00000000";
		ram_buffer(8094) := X"00000000";
		ram_buffer(8095) := X"00000000";
		ram_buffer(8096) := X"00000000";
		ram_buffer(8097) := X"00000000";
		ram_buffer(8098) := X"00000000";
		ram_buffer(8099) := X"00000000";
		ram_buffer(8100) := X"00000000";
		ram_buffer(8101) := X"00000000";
		ram_buffer(8102) := X"00000000";
		ram_buffer(8103) := X"00000000";
		ram_buffer(8104) := X"00000000";
		ram_buffer(8105) := X"00000000";
		ram_buffer(8106) := X"00000000";
		ram_buffer(8107) := X"00000000";
		ram_buffer(8108) := X"00000000";
		ram_buffer(8109) := X"00000000";
		ram_buffer(8110) := X"00000000";
		ram_buffer(8111) := X"00000000";
		ram_buffer(8112) := X"00000000";
		ram_buffer(8113) := X"00000000";
		ram_buffer(8114) := X"00000000";
		ram_buffer(8115) := X"00000000";
		ram_buffer(8116) := X"00000000";
		ram_buffer(8117) := X"00000000";
		ram_buffer(8118) := X"00000000";
		ram_buffer(8119) := X"00000000";
		ram_buffer(8120) := X"00000000";
		ram_buffer(8121) := X"00000000";
		ram_buffer(8122) := X"00000000";
		ram_buffer(8123) := X"00000000";
		ram_buffer(8124) := X"00000000";
		ram_buffer(8125) := X"00000000";
		ram_buffer(8126) := X"00000000";
		ram_buffer(8127) := X"00000000";
		ram_buffer(8128) := X"00000000";
		ram_buffer(8129) := X"00000000";
		ram_buffer(8130) := X"00000000";
		ram_buffer(8131) := X"00000000";
		ram_buffer(8132) := X"00000000";
		ram_buffer(8133) := X"00000000";
		ram_buffer(8134) := X"00000000";
		ram_buffer(8135) := X"00000000";
		ram_buffer(8136) := X"00000000";
		ram_buffer(8137) := X"00000000";
		ram_buffer(8138) := X"00000000";
		ram_buffer(8139) := X"00000000";
		ram_buffer(8140) := X"00000000";
		ram_buffer(8141) := X"00000000";
		ram_buffer(8142) := X"00000000";
		ram_buffer(8143) := X"00000000";
		ram_buffer(8144) := X"00000000";
		ram_buffer(8145) := X"00000000";
		ram_buffer(8146) := X"00000000";
		ram_buffer(8147) := X"00000000";
		ram_buffer(8148) := X"00000000";
		ram_buffer(8149) := X"00000000";
		ram_buffer(8150) := X"00000000";
		ram_buffer(8151) := X"00000000";
		ram_buffer(8152) := X"00000000";
		ram_buffer(8153) := X"00000000";
		ram_buffer(8154) := X"00000000";
		ram_buffer(8155) := X"00000000";
		ram_buffer(8156) := X"00000000";
		ram_buffer(8157) := X"00000000";
		ram_buffer(8158) := X"00000000";
		ram_buffer(8159) := X"00000000";
		ram_buffer(8160) := X"00000000";
		ram_buffer(8161) := X"00000000";
		ram_buffer(8162) := X"00000000";
		ram_buffer(8163) := X"00000000";
		ram_buffer(8164) := X"00000000";
		ram_buffer(8165) := X"00000000";
		ram_buffer(8166) := X"00000000";
		ram_buffer(8167) := X"00000000";
		ram_buffer(8168) := X"00000000";
		ram_buffer(8169) := X"00000000";
		ram_buffer(8170) := X"00000000";
		ram_buffer(8171) := X"00000000";
		ram_buffer(8172) := X"00000000";
		ram_buffer(8173) := X"00000000";
		ram_buffer(8174) := X"00000000";
		ram_buffer(8175) := X"00000000";
		ram_buffer(8176) := X"00000000";
		ram_buffer(8177) := X"00000000";
		ram_buffer(8178) := X"00000000";
		ram_buffer(8179) := X"00000000";
		ram_buffer(8180) := X"00000000";
		ram_buffer(8181) := X"00000000";
		ram_buffer(8182) := X"00000000";
		ram_buffer(8183) := X"00000000";
		ram_buffer(8184) := X"00000000";
		ram_buffer(8185) := X"00000000";
		ram_buffer(8186) := X"00000000";
		ram_buffer(8187) := X"00000000";
		ram_buffer(8188) := X"00000000";
		ram_buffer(8189) := X"00000000";
		ram_buffer(8190) := X"00000000";
		ram_buffer(8191) := X"00000000";
		ram_buffer(8192) := X"00000000";
		ram_buffer(8193) := X"00000000";
		ram_buffer(8194) := X"00000000";
		ram_buffer(8195) := X"00000000";
		ram_buffer(8196) := X"00000000";
		ram_buffer(8197) := X"00000000";
		ram_buffer(8198) := X"00000000";
		ram_buffer(8199) := X"00000000";
		ram_buffer(8200) := X"00000000";
		ram_buffer(8201) := X"00000000";
		ram_buffer(8202) := X"00000000";
		ram_buffer(8203) := X"00000000";
		ram_buffer(8204) := X"00000000";
		ram_buffer(8205) := X"00000000";
		ram_buffer(8206) := X"00000000";
		ram_buffer(8207) := X"00000000";
		ram_buffer(8208) := X"00000000";
		ram_buffer(8209) := X"00000000";
		ram_buffer(8210) := X"00000000";
		ram_buffer(8211) := X"00000000";
		ram_buffer(8212) := X"00000000";
		ram_buffer(8213) := X"00000000";
		ram_buffer(8214) := X"00000000";
		ram_buffer(8215) := X"00000000";
		ram_buffer(8216) := X"00000000";
		ram_buffer(8217) := X"00000000";
		ram_buffer(8218) := X"00000000";
		ram_buffer(8219) := X"00000000";
		ram_buffer(8220) := X"00000000";
		ram_buffer(8221) := X"00000000";
		ram_buffer(8222) := X"00000000";
		ram_buffer(8223) := X"00000000";
		ram_buffer(8224) := X"00000000";
		ram_buffer(8225) := X"00000000";
		ram_buffer(8226) := X"00000000";
		ram_buffer(8227) := X"00000000";
		ram_buffer(8228) := X"00000000";
		ram_buffer(8229) := X"00000000";
		ram_buffer(8230) := X"00000000";
		ram_buffer(8231) := X"00000000";
		ram_buffer(8232) := X"00000000";
		ram_buffer(8233) := X"00000000";
		ram_buffer(8234) := X"00000000";
		ram_buffer(8235) := X"00000000";
		ram_buffer(8236) := X"00000000";
		ram_buffer(8237) := X"00000000";
		ram_buffer(8238) := X"00000000";
		ram_buffer(8239) := X"00000000";
		ram_buffer(8240) := X"00000000";
		ram_buffer(8241) := X"00000000";
		ram_buffer(8242) := X"00000000";
		ram_buffer(8243) := X"00000000";
		ram_buffer(8244) := X"00000000";
		ram_buffer(8245) := X"00000000";
		ram_buffer(8246) := X"00000000";
		ram_buffer(8247) := X"00000000";
		ram_buffer(8248) := X"00000000";
		ram_buffer(8249) := X"00000000";
		ram_buffer(8250) := X"00000000";
		ram_buffer(8251) := X"00000000";
		ram_buffer(8252) := X"00000000";
		ram_buffer(8253) := X"00000000";
		ram_buffer(8254) := X"00000000";
		ram_buffer(8255) := X"00000000";
		ram_buffer(8256) := X"00000000";
		ram_buffer(8257) := X"00000000";
		ram_buffer(8258) := X"00000000";
		ram_buffer(8259) := X"00000000";
		ram_buffer(8260) := X"00000000";
		ram_buffer(8261) := X"00000000";
		ram_buffer(8262) := X"00000000";
		ram_buffer(8263) := X"00000000";
		ram_buffer(8264) := X"00000000";
		ram_buffer(8265) := X"00000000";
		ram_buffer(8266) := X"00000000";
		ram_buffer(8267) := X"00000000";
		ram_buffer(8268) := X"00000000";
		ram_buffer(8269) := X"00000000";
		ram_buffer(8270) := X"00000000";
		ram_buffer(8271) := X"00000000";
		ram_buffer(8272) := X"00000000";
		ram_buffer(8273) := X"00000000";
		ram_buffer(8274) := X"00000000";
		ram_buffer(8275) := X"00000000";
		ram_buffer(8276) := X"00000000";
		ram_buffer(8277) := X"00000000";
		ram_buffer(8278) := X"00000000";
		ram_buffer(8279) := X"00000000";
		ram_buffer(8280) := X"00000000";
		ram_buffer(8281) := X"00000000";
		ram_buffer(8282) := X"00000000";
		ram_buffer(8283) := X"00000000";
		ram_buffer(8284) := X"00000000";
		ram_buffer(8285) := X"00000000";
		ram_buffer(8286) := X"00000000";
		ram_buffer(8287) := X"00000000";
		ram_buffer(8288) := X"00000000";
		ram_buffer(8289) := X"00000000";
		ram_buffer(8290) := X"00000000";
		ram_buffer(8291) := X"00000000";
		ram_buffer(8292) := X"00000000";
		ram_buffer(8293) := X"00000000";
		ram_buffer(8294) := X"00000000";
		ram_buffer(8295) := X"00000000";
		ram_buffer(8296) := X"00000000";
		ram_buffer(8297) := X"00000000";
		ram_buffer(8298) := X"00000000";
		ram_buffer(8299) := X"00000000";
		ram_buffer(8300) := X"00000000";
		ram_buffer(8301) := X"00000000";
		ram_buffer(8302) := X"00000000";
		ram_buffer(8303) := X"00000000";
		ram_buffer(8304) := X"00000000";
		ram_buffer(8305) := X"00000000";
		ram_buffer(8306) := X"00000000";
		ram_buffer(8307) := X"00000000";
		ram_buffer(8308) := X"00000000";
		ram_buffer(8309) := X"00000000";
		ram_buffer(8310) := X"00000000";
		ram_buffer(8311) := X"00000000";
		ram_buffer(8312) := X"00000000";
		ram_buffer(8313) := X"00000000";
		ram_buffer(8314) := X"00000000";
		ram_buffer(8315) := X"00000000";
		ram_buffer(8316) := X"00000000";
		ram_buffer(8317) := X"00000000";
		ram_buffer(8318) := X"00000000";
		ram_buffer(8319) := X"00000000";
		ram_buffer(8320) := X"00000000";
		ram_buffer(8321) := X"00000000";
		ram_buffer(8322) := X"00000000";
		ram_buffer(8323) := X"00000000";
		ram_buffer(8324) := X"00000000";
		ram_buffer(8325) := X"00000000";
		ram_buffer(8326) := X"00000000";
		ram_buffer(8327) := X"00000000";
		ram_buffer(8328) := X"00000000";
		ram_buffer(8329) := X"00000000";
		ram_buffer(8330) := X"00000000";
		ram_buffer(8331) := X"00000000";
		ram_buffer(8332) := X"00000000";
		ram_buffer(8333) := X"00000000";
		ram_buffer(8334) := X"00000000";
		ram_buffer(8335) := X"00000000";
		ram_buffer(8336) := X"00000000";
		ram_buffer(8337) := X"00000000";
		ram_buffer(8338) := X"00000000";
		ram_buffer(8339) := X"00000000";
		ram_buffer(8340) := X"00000000";
		ram_buffer(8341) := X"00000000";
		ram_buffer(8342) := X"00000000";
		ram_buffer(8343) := X"00000000";
		ram_buffer(8344) := X"00000000";
		ram_buffer(8345) := X"00000000";
		ram_buffer(8346) := X"00000000";
		ram_buffer(8347) := X"00000000";
		ram_buffer(8348) := X"00000000";
		ram_buffer(8349) := X"00000000";
		ram_buffer(8350) := X"00000000";
		ram_buffer(8351) := X"00000000";
		ram_buffer(8352) := X"00000000";
		ram_buffer(8353) := X"00000000";
		ram_buffer(8354) := X"00000000";
		ram_buffer(8355) := X"00000000";
		ram_buffer(8356) := X"00000000";
		ram_buffer(8357) := X"00000000";
		ram_buffer(8358) := X"00000000";
		ram_buffer(8359) := X"00000000";
		ram_buffer(8360) := X"00000000";
		ram_buffer(8361) := X"00000000";
		ram_buffer(8362) := X"00000000";
		ram_buffer(8363) := X"00000000";
		ram_buffer(8364) := X"00000000";
		ram_buffer(8365) := X"00000000";
		ram_buffer(8366) := X"00000000";
		ram_buffer(8367) := X"00000000";
		ram_buffer(8368) := X"00000000";
		ram_buffer(8369) := X"00000000";
		ram_buffer(8370) := X"00000000";
		ram_buffer(8371) := X"00000000";
		ram_buffer(8372) := X"00000000";
		ram_buffer(8373) := X"00000000";
		ram_buffer(8374) := X"00000000";
		ram_buffer(8375) := X"00000000";
		ram_buffer(8376) := X"00000000";
		ram_buffer(8377) := X"00000000";
		ram_buffer(8378) := X"00000000";
		ram_buffer(8379) := X"00000000";
		ram_buffer(8380) := X"00000000";
		ram_buffer(8381) := X"00000000";
		ram_buffer(8382) := X"00000000";
		ram_buffer(8383) := X"00000000";
		ram_buffer(8384) := X"00000000";
		ram_buffer(8385) := X"00000000";
		ram_buffer(8386) := X"00000000";
		ram_buffer(8387) := X"00000000";
		ram_buffer(8388) := X"00000000";
		ram_buffer(8389) := X"00000000";
		ram_buffer(8390) := X"00000000";
		ram_buffer(8391) := X"00000000";
		ram_buffer(8392) := X"00000000";
		ram_buffer(8393) := X"00000000";
		ram_buffer(8394) := X"00000000";
		ram_buffer(8395) := X"00000000";
		ram_buffer(8396) := X"00000000";
		ram_buffer(8397) := X"00000000";
		ram_buffer(8398) := X"00000000";
		ram_buffer(8399) := X"00000000";
		ram_buffer(8400) := X"00000000";
		ram_buffer(8401) := X"00000000";
		ram_buffer(8402) := X"00000000";
		ram_buffer(8403) := X"00000000";
		ram_buffer(8404) := X"00000000";
		ram_buffer(8405) := X"00000000";
		ram_buffer(8406) := X"00000000";
		ram_buffer(8407) := X"00000000";
		ram_buffer(8408) := X"00000000";
		ram_buffer(8409) := X"00000000";
		ram_buffer(8410) := X"00000000";
		ram_buffer(8411) := X"00000000";
		ram_buffer(8412) := X"00000000";
		ram_buffer(8413) := X"00000000";
		ram_buffer(8414) := X"00000000";
		ram_buffer(8415) := X"00000000";
		ram_buffer(8416) := X"00000000";
		ram_buffer(8417) := X"00000000";
		ram_buffer(8418) := X"00000000";
		ram_buffer(8419) := X"00000000";
		ram_buffer(8420) := X"00000000";
		ram_buffer(8421) := X"00000000";
		ram_buffer(8422) := X"00000000";
		ram_buffer(8423) := X"00000000";
		ram_buffer(8424) := X"00000000";
		ram_buffer(8425) := X"00000000";
		ram_buffer(8426) := X"00000000";
		ram_buffer(8427) := X"00000000";
		ram_buffer(8428) := X"00000000";
		ram_buffer(8429) := X"00000000";
		ram_buffer(8430) := X"00000000";
		ram_buffer(8431) := X"00000000";
		ram_buffer(8432) := X"00000000";
		ram_buffer(8433) := X"00000000";
		ram_buffer(8434) := X"00000000";
		ram_buffer(8435) := X"00000000";
		ram_buffer(8436) := X"00000000";
		ram_buffer(8437) := X"00000000";
		ram_buffer(8438) := X"00000000";
		ram_buffer(8439) := X"00000000";
		ram_buffer(8440) := X"00000000";
		ram_buffer(8441) := X"00000000";
		ram_buffer(8442) := X"00000000";
		ram_buffer(8443) := X"00000000";
		ram_buffer(8444) := X"00000000";
		ram_buffer(8445) := X"00000000";
		ram_buffer(8446) := X"00000000";
		ram_buffer(8447) := X"00000000";
		ram_buffer(8448) := X"00000000";
		ram_buffer(8449) := X"00000000";
		ram_buffer(8450) := X"00000000";
		ram_buffer(8451) := X"00000000";
		ram_buffer(8452) := X"00000000";
		ram_buffer(8453) := X"00000000";
		ram_buffer(8454) := X"00000000";
		ram_buffer(8455) := X"00000000";
		ram_buffer(8456) := X"00000000";
		ram_buffer(8457) := X"00000000";
		ram_buffer(8458) := X"00000000";
		ram_buffer(8459) := X"00000000";
		ram_buffer(8460) := X"00000000";
		ram_buffer(8461) := X"00000000";
		ram_buffer(8462) := X"00000000";
		ram_buffer(8463) := X"00000000";
		ram_buffer(8464) := X"00000000";
		ram_buffer(8465) := X"00000000";
		ram_buffer(8466) := X"00000000";
		ram_buffer(8467) := X"00000000";
		ram_buffer(8468) := X"00000000";
		ram_buffer(8469) := X"00000000";
		ram_buffer(8470) := X"00000000";
		ram_buffer(8471) := X"00000000";
		ram_buffer(8472) := X"00000000";
		ram_buffer(8473) := X"00000000";
		ram_buffer(8474) := X"00000000";
		ram_buffer(8475) := X"00000000";
		ram_buffer(8476) := X"00000000";
		ram_buffer(8477) := X"00000000";
		ram_buffer(8478) := X"00000000";
		ram_buffer(8479) := X"00000000";
		ram_buffer(8480) := X"00000000";
		ram_buffer(8481) := X"00000000";
		ram_buffer(8482) := X"00000000";
		ram_buffer(8483) := X"00000000";
		ram_buffer(8484) := X"00000000";
		ram_buffer(8485) := X"00000000";
		ram_buffer(8486) := X"00000000";
		ram_buffer(8487) := X"00000000";
		ram_buffer(8488) := X"00000000";
		ram_buffer(8489) := X"00000000";
		ram_buffer(8490) := X"00000000";
		ram_buffer(8491) := X"00000000";
		ram_buffer(8492) := X"00000000";
		ram_buffer(8493) := X"00000000";
		ram_buffer(8494) := X"00000000";
		ram_buffer(8495) := X"00000000";
		ram_buffer(8496) := X"00000000";
		ram_buffer(8497) := X"00000000";
		ram_buffer(8498) := X"00000000";
		ram_buffer(8499) := X"00000000";
		ram_buffer(8500) := X"00000000";
		ram_buffer(8501) := X"00000000";
		ram_buffer(8502) := X"00000000";
		ram_buffer(8503) := X"00000000";
		ram_buffer(8504) := X"00000000";
		ram_buffer(8505) := X"00000000";
		ram_buffer(8506) := X"00000000";
		ram_buffer(8507) := X"00000000";
		ram_buffer(8508) := X"00000000";
		ram_buffer(8509) := X"00000000";
		ram_buffer(8510) := X"00000000";
		ram_buffer(8511) := X"00000000";
		ram_buffer(8512) := X"00000000";
		ram_buffer(8513) := X"00000000";
		ram_buffer(8514) := X"00000000";
		ram_buffer(8515) := X"00000000";
		ram_buffer(8516) := X"00000000";
		ram_buffer(8517) := X"00000000";
		ram_buffer(8518) := X"00000000";
		ram_buffer(8519) := X"00000000";
		ram_buffer(8520) := X"00000000";
		ram_buffer(8521) := X"00000000";
		ram_buffer(8522) := X"00000000";
		ram_buffer(8523) := X"00000000";
		ram_buffer(8524) := X"00000000";
		ram_buffer(8525) := X"00000000";
		ram_buffer(8526) := X"00000000";
		ram_buffer(8527) := X"00000000";
		ram_buffer(8528) := X"00000000";
		ram_buffer(8529) := X"00000000";
		ram_buffer(8530) := X"00000000";
		ram_buffer(8531) := X"00000000";
		ram_buffer(8532) := X"00000000";
		ram_buffer(8533) := X"00000000";
		ram_buffer(8534) := X"00000000";
		ram_buffer(8535) := X"00000000";
		ram_buffer(8536) := X"00000000";
		ram_buffer(8537) := X"00000000";
		ram_buffer(8538) := X"00000000";
		ram_buffer(8539) := X"00000000";
		ram_buffer(8540) := X"00000000";
		ram_buffer(8541) := X"00000000";
		ram_buffer(8542) := X"00000000";
		ram_buffer(8543) := X"00000000";
		ram_buffer(8544) := X"00000000";
		ram_buffer(8545) := X"00000000";
		ram_buffer(8546) := X"00000000";
		ram_buffer(8547) := X"00000000";
		ram_buffer(8548) := X"00000000";
		ram_buffer(8549) := X"00000000";
		ram_buffer(8550) := X"00000000";
		ram_buffer(8551) := X"00000000";
		ram_buffer(8552) := X"00000000";
		ram_buffer(8553) := X"00000000";
		ram_buffer(8554) := X"00000000";
		ram_buffer(8555) := X"00000000";
		ram_buffer(8556) := X"00000000";
		ram_buffer(8557) := X"00000000";
		ram_buffer(8558) := X"00000000";
		ram_buffer(8559) := X"00000000";
		ram_buffer(8560) := X"00000000";
		ram_buffer(8561) := X"00000000";
		ram_buffer(8562) := X"00000000";
		ram_buffer(8563) := X"00000000";
		ram_buffer(8564) := X"00000000";
		ram_buffer(8565) := X"00000000";
		ram_buffer(8566) := X"00000000";
		ram_buffer(8567) := X"00000000";
		ram_buffer(8568) := X"00000000";
		ram_buffer(8569) := X"00000000";
		ram_buffer(8570) := X"00000000";
		ram_buffer(8571) := X"00000000";
		ram_buffer(8572) := X"00000000";
		ram_buffer(8573) := X"00000000";
		ram_buffer(8574) := X"00000000";
		ram_buffer(8575) := X"00000000";
		ram_buffer(8576) := X"00000000";
		ram_buffer(8577) := X"00000000";
		ram_buffer(8578) := X"00000000";
		ram_buffer(8579) := X"00000000";
		ram_buffer(8580) := X"00000000";
		ram_buffer(8581) := X"00000000";
		ram_buffer(8582) := X"00000000";
		ram_buffer(8583) := X"00000000";
		ram_buffer(8584) := X"00000000";
		ram_buffer(8585) := X"00000000";
		ram_buffer(8586) := X"00000000";
		ram_buffer(8587) := X"00000000";
		ram_buffer(8588) := X"00000000";
		ram_buffer(8589) := X"00000000";
		ram_buffer(8590) := X"00000000";
		ram_buffer(8591) := X"00000000";
		ram_buffer(8592) := X"00000000";
		ram_buffer(8593) := X"00000000";
		ram_buffer(8594) := X"00000000";
		ram_buffer(8595) := X"00000000";
		ram_buffer(8596) := X"00000000";
		ram_buffer(8597) := X"00000000";
		ram_buffer(8598) := X"00000000";
		ram_buffer(8599) := X"00000000";
		ram_buffer(8600) := X"00000000";
		ram_buffer(8601) := X"00000000";
		ram_buffer(8602) := X"00000000";
		ram_buffer(8603) := X"00000000";
		ram_buffer(8604) := X"00000000";
		ram_buffer(8605) := X"00000000";
		ram_buffer(8606) := X"00000000";
		ram_buffer(8607) := X"00000000";
		ram_buffer(8608) := X"00000000";
		ram_buffer(8609) := X"00000000";
		ram_buffer(8610) := X"00000000";
		ram_buffer(8611) := X"00000000";
		ram_buffer(8612) := X"00000000";
		ram_buffer(8613) := X"00000000";
		ram_buffer(8614) := X"00000000";
		ram_buffer(8615) := X"00000000";
		ram_buffer(8616) := X"00000000";
		ram_buffer(8617) := X"00000000";
		ram_buffer(8618) := X"00000000";
		ram_buffer(8619) := X"00000000";
		ram_buffer(8620) := X"00000000";
		ram_buffer(8621) := X"00000000";
		ram_buffer(8622) := X"00000000";
		ram_buffer(8623) := X"00000000";
		ram_buffer(8624) := X"00000000";
		ram_buffer(8625) := X"00000000";
		ram_buffer(8626) := X"00000000";
		ram_buffer(8627) := X"00000000";
		ram_buffer(8628) := X"00000000";
		ram_buffer(8629) := X"00000000";
		ram_buffer(8630) := X"00000000";
		ram_buffer(8631) := X"00000000";
		ram_buffer(8632) := X"00000000";
		ram_buffer(8633) := X"00000000";
		ram_buffer(8634) := X"00000000";
		ram_buffer(8635) := X"00000000";
		ram_buffer(8636) := X"00000000";
		ram_buffer(8637) := X"00000000";
		ram_buffer(8638) := X"00000000";
		ram_buffer(8639) := X"00000000";
		ram_buffer(8640) := X"00000000";
		ram_buffer(8641) := X"00000000";
		ram_buffer(8642) := X"00000000";
		ram_buffer(8643) := X"00000000";
		ram_buffer(8644) := X"00000000";
		ram_buffer(8645) := X"00000000";
		ram_buffer(8646) := X"00000000";
		ram_buffer(8647) := X"00000000";
		ram_buffer(8648) := X"00000000";
		ram_buffer(8649) := X"00000000";
		ram_buffer(8650) := X"00000000";
		ram_buffer(8651) := X"00000000";
		ram_buffer(8652) := X"00000000";
		ram_buffer(8653) := X"00000000";
		ram_buffer(8654) := X"00000000";
		ram_buffer(8655) := X"00000000";
		ram_buffer(8656) := X"00000000";
		ram_buffer(8657) := X"00000000";
		ram_buffer(8658) := X"00000000";
		ram_buffer(8659) := X"00000000";
		ram_buffer(8660) := X"00000000";
		ram_buffer(8661) := X"00000000";
		ram_buffer(8662) := X"00000000";
		ram_buffer(8663) := X"00000000";
		ram_buffer(8664) := X"00000000";
		ram_buffer(8665) := X"00000000";
		ram_buffer(8666) := X"00000000";
		ram_buffer(8667) := X"00000000";
		ram_buffer(8668) := X"00000000";
		ram_buffer(8669) := X"00000000";
		ram_buffer(8670) := X"00000000";
		ram_buffer(8671) := X"00000000";
		ram_buffer(8672) := X"00000000";
		ram_buffer(8673) := X"00000000";
		ram_buffer(8674) := X"00000000";
		ram_buffer(8675) := X"00000000";
		ram_buffer(8676) := X"00000000";
		ram_buffer(8677) := X"00000000";
		ram_buffer(8678) := X"00000000";
		ram_buffer(8679) := X"00000000";
		ram_buffer(8680) := X"00000000";
		ram_buffer(8681) := X"00000000";
		ram_buffer(8682) := X"00000000";
		ram_buffer(8683) := X"00000000";
		ram_buffer(8684) := X"00000000";
		ram_buffer(8685) := X"00000000";
		ram_buffer(8686) := X"00000000";
		ram_buffer(8687) := X"00000000";
		ram_buffer(8688) := X"00000000";
		ram_buffer(8689) := X"00000000";
		ram_buffer(8690) := X"00000000";
		ram_buffer(8691) := X"00000000";
		ram_buffer(8692) := X"00000000";
		ram_buffer(8693) := X"00000000";
		ram_buffer(8694) := X"00000000";
		ram_buffer(8695) := X"00000000";
		ram_buffer(8696) := X"00000000";
		ram_buffer(8697) := X"00000000";
		ram_buffer(8698) := X"00000000";
		ram_buffer(8699) := X"00000000";
		ram_buffer(8700) := X"00000000";
		ram_buffer(8701) := X"00000000";
		ram_buffer(8702) := X"00000000";
		ram_buffer(8703) := X"00000000";
		ram_buffer(8704) := X"00000000";
		ram_buffer(8705) := X"00000000";
		ram_buffer(8706) := X"00000000";
		ram_buffer(8707) := X"00000000";
		ram_buffer(8708) := X"00000000";
		ram_buffer(8709) := X"00000000";
		ram_buffer(8710) := X"00000000";
		ram_buffer(8711) := X"00000000";
		ram_buffer(8712) := X"00000000";
		ram_buffer(8713) := X"00000000";
		ram_buffer(8714) := X"00000000";
		ram_buffer(8715) := X"00000000";
		ram_buffer(8716) := X"00000000";
		ram_buffer(8717) := X"00000000";
		ram_buffer(8718) := X"00000000";
		ram_buffer(8719) := X"00000000";
		ram_buffer(8720) := X"00000000";
		ram_buffer(8721) := X"00000000";
		ram_buffer(8722) := X"00000000";
		ram_buffer(8723) := X"00000000";
		ram_buffer(8724) := X"00000000";
		ram_buffer(8725) := X"00000000";
		ram_buffer(8726) := X"00000000";
		ram_buffer(8727) := X"00000000";
		ram_buffer(8728) := X"00000000";
		ram_buffer(8729) := X"00000000";
		ram_buffer(8730) := X"00000000";
		ram_buffer(8731) := X"00000000";
		ram_buffer(8732) := X"00000000";
		ram_buffer(8733) := X"00000000";
		ram_buffer(8734) := X"00000000";
		ram_buffer(8735) := X"00000000";
		ram_buffer(8736) := X"00000000";
		ram_buffer(8737) := X"00000000";
		ram_buffer(8738) := X"00000000";
		ram_buffer(8739) := X"00000000";
		ram_buffer(8740) := X"00000000";
		ram_buffer(8741) := X"00000000";
		ram_buffer(8742) := X"00000000";
		ram_buffer(8743) := X"00000000";
		ram_buffer(8744) := X"00000000";
		ram_buffer(8745) := X"00000000";
		ram_buffer(8746) := X"00000000";
		ram_buffer(8747) := X"00000000";
		ram_buffer(8748) := X"00000000";
		ram_buffer(8749) := X"00000000";
		ram_buffer(8750) := X"00000000";
		ram_buffer(8751) := X"00000000";
		ram_buffer(8752) := X"00000000";
		ram_buffer(8753) := X"00000000";
		ram_buffer(8754) := X"00000000";
		ram_buffer(8755) := X"00000000";
		ram_buffer(8756) := X"00000000";
		ram_buffer(8757) := X"00000000";
		ram_buffer(8758) := X"00000000";
		ram_buffer(8759) := X"00000000";
		ram_buffer(8760) := X"00000000";
		ram_buffer(8761) := X"00000000";
		ram_buffer(8762) := X"00000000";
		ram_buffer(8763) := X"00000000";
		ram_buffer(8764) := X"00000000";
		ram_buffer(8765) := X"00000000";
		ram_buffer(8766) := X"00000000";
		ram_buffer(8767) := X"00000000";
		ram_buffer(8768) := X"00000000";
		ram_buffer(8769) := X"00000000";
		ram_buffer(8770) := X"00000000";
		ram_buffer(8771) := X"00000000";
		ram_buffer(8772) := X"00000000";
		ram_buffer(8773) := X"00000000";
		ram_buffer(8774) := X"00000000";
		ram_buffer(8775) := X"00000000";
		ram_buffer(8776) := X"00000000";
		ram_buffer(8777) := X"00000000";
		ram_buffer(8778) := X"00000000";
		ram_buffer(8779) := X"00000000";
		ram_buffer(8780) := X"00000000";
		ram_buffer(8781) := X"00000000";
		ram_buffer(8782) := X"00000000";
		ram_buffer(8783) := X"00000000";
		ram_buffer(8784) := X"00000000";
		ram_buffer(8785) := X"00000000";
		ram_buffer(8786) := X"00000000";
		ram_buffer(8787) := X"00000000";
		ram_buffer(8788) := X"00000000";
		ram_buffer(8789) := X"00000000";
		ram_buffer(8790) := X"00000000";
		ram_buffer(8791) := X"00000000";
		ram_buffer(8792) := X"00000000";
		ram_buffer(8793) := X"00000000";
		ram_buffer(8794) := X"00000000";
		ram_buffer(8795) := X"00000000";
		ram_buffer(8796) := X"00000000";
		ram_buffer(8797) := X"00000000";
		ram_buffer(8798) := X"00000000";
		ram_buffer(8799) := X"00000000";
		ram_buffer(8800) := X"00000000";
		ram_buffer(8801) := X"00000000";
		ram_buffer(8802) := X"00000000";
		ram_buffer(8803) := X"00000000";
		ram_buffer(8804) := X"00000000";
		ram_buffer(8805) := X"00000000";
		ram_buffer(8806) := X"00000000";
		ram_buffer(8807) := X"00000000";
		ram_buffer(8808) := X"00000000";
		ram_buffer(8809) := X"00000000";
		ram_buffer(8810) := X"00000000";
		ram_buffer(8811) := X"00000000";
		ram_buffer(8812) := X"00000000";
		ram_buffer(8813) := X"00000000";
		ram_buffer(8814) := X"00000000";
		ram_buffer(8815) := X"00000000";
		ram_buffer(8816) := X"00000000";
		ram_buffer(8817) := X"00000000";
		ram_buffer(8818) := X"00000000";
		ram_buffer(8819) := X"00000000";
		ram_buffer(8820) := X"00000000";
		ram_buffer(8821) := X"00000000";
		ram_buffer(8822) := X"00000000";
		ram_buffer(8823) := X"00000000";
		ram_buffer(8824) := X"00000000";
		ram_buffer(8825) := X"00000000";
		ram_buffer(8826) := X"00000000";
		ram_buffer(8827) := X"00000000";
		ram_buffer(8828) := X"00000000";
		ram_buffer(8829) := X"00000000";
		ram_buffer(8830) := X"00000000";
		ram_buffer(8831) := X"00000000";
		ram_buffer(8832) := X"00000000";
		ram_buffer(8833) := X"00000000";
		ram_buffer(8834) := X"00000000";
		ram_buffer(8835) := X"00000000";
		ram_buffer(8836) := X"00000000";
		ram_buffer(8837) := X"00000000";
		ram_buffer(8838) := X"00000000";
		ram_buffer(8839) := X"00000000";
		ram_buffer(8840) := X"00000000";
		ram_buffer(8841) := X"00000000";
		ram_buffer(8842) := X"00000000";
		ram_buffer(8843) := X"00000000";
		ram_buffer(8844) := X"00000000";
		ram_buffer(8845) := X"00000000";
		ram_buffer(8846) := X"00000000";
		ram_buffer(8847) := X"00000000";
		ram_buffer(8848) := X"00000000";
		ram_buffer(8849) := X"00000000";
		ram_buffer(8850) := X"00000000";
		ram_buffer(8851) := X"00000000";
		ram_buffer(8852) := X"00000000";
		ram_buffer(8853) := X"00000000";
		ram_buffer(8854) := X"00000000";
		ram_buffer(8855) := X"00000000";
		ram_buffer(8856) := X"00000000";
		ram_buffer(8857) := X"00000000";
		ram_buffer(8858) := X"00000000";
		ram_buffer(8859) := X"00000000";
		ram_buffer(8860) := X"00000000";
		ram_buffer(8861) := X"00000000";
		ram_buffer(8862) := X"00000000";
		ram_buffer(8863) := X"00000000";
		ram_buffer(8864) := X"00000000";
		ram_buffer(8865) := X"00000000";
		ram_buffer(8866) := X"00000000";
		ram_buffer(8867) := X"00000000";
		ram_buffer(8868) := X"00000000";
		ram_buffer(8869) := X"00000000";
		ram_buffer(8870) := X"00000000";
		ram_buffer(8871) := X"00000000";
		ram_buffer(8872) := X"00000000";
		ram_buffer(8873) := X"00000000";
		ram_buffer(8874) := X"00000000";
		ram_buffer(8875) := X"00000000";
		ram_buffer(8876) := X"00000000";
		ram_buffer(8877) := X"00000000";
		ram_buffer(8878) := X"00000000";
		ram_buffer(8879) := X"00000000";
		ram_buffer(8880) := X"00000000";
		ram_buffer(8881) := X"00000000";
		ram_buffer(8882) := X"00000000";
		ram_buffer(8883) := X"00000000";
		ram_buffer(8884) := X"00000000";
		ram_buffer(8885) := X"00000000";
		ram_buffer(8886) := X"00000000";
		ram_buffer(8887) := X"00000000";
		ram_buffer(8888) := X"00000000";
		ram_buffer(8889) := X"00000000";
		ram_buffer(8890) := X"00000000";
		ram_buffer(8891) := X"00000000";
		ram_buffer(8892) := X"00000000";
		ram_buffer(8893) := X"00000000";
		ram_buffer(8894) := X"00000000";
		ram_buffer(8895) := X"00000000";
		ram_buffer(8896) := X"00000000";
		ram_buffer(8897) := X"00000000";
		ram_buffer(8898) := X"00000000";
		ram_buffer(8899) := X"00000000";
		ram_buffer(8900) := X"00000000";
		ram_buffer(8901) := X"00000000";
		ram_buffer(8902) := X"00000000";
		ram_buffer(8903) := X"00000000";
		ram_buffer(8904) := X"00000000";
		ram_buffer(8905) := X"00000000";
		ram_buffer(8906) := X"00000000";
		ram_buffer(8907) := X"00000000";
		ram_buffer(8908) := X"00000000";
		ram_buffer(8909) := X"00000000";
		ram_buffer(8910) := X"00000000";
		ram_buffer(8911) := X"00000000";
		ram_buffer(8912) := X"00000000";
		ram_buffer(8913) := X"00000000";
		ram_buffer(8914) := X"00000000";
		ram_buffer(8915) := X"00000000";
		ram_buffer(8916) := X"00000000";
		ram_buffer(8917) := X"00000000";
		ram_buffer(8918) := X"00000000";
		ram_buffer(8919) := X"00000000";
		ram_buffer(8920) := X"00000000";
		ram_buffer(8921) := X"00000000";
		ram_buffer(8922) := X"00000000";
		ram_buffer(8923) := X"00000000";
		ram_buffer(8924) := X"00000000";
		ram_buffer(8925) := X"00000000";
		ram_buffer(8926) := X"00000000";
		ram_buffer(8927) := X"00000000";
		ram_buffer(8928) := X"00000000";
		ram_buffer(8929) := X"00000000";
		ram_buffer(8930) := X"00000000";
		ram_buffer(8931) := X"00000000";
		ram_buffer(8932) := X"00000000";
		ram_buffer(8933) := X"00000000";
		ram_buffer(8934) := X"00000000";
		ram_buffer(8935) := X"00000000";
		ram_buffer(8936) := X"00000000";
		ram_buffer(8937) := X"00000000";
		ram_buffer(8938) := X"00000000";
		ram_buffer(8939) := X"00000000";
		ram_buffer(8940) := X"00000000";
		ram_buffer(8941) := X"00000000";
		ram_buffer(8942) := X"00000000";
		ram_buffer(8943) := X"00000000";
		ram_buffer(8944) := X"00000000";
		ram_buffer(8945) := X"00000000";
		ram_buffer(8946) := X"00000000";
		ram_buffer(8947) := X"00000000";
		ram_buffer(8948) := X"00000000";
		ram_buffer(8949) := X"00000000";
		ram_buffer(8950) := X"00000000";
		ram_buffer(8951) := X"00000000";
		ram_buffer(8952) := X"00000000";
		ram_buffer(8953) := X"00000000";
		ram_buffer(8954) := X"00000000";
		ram_buffer(8955) := X"00000000";
		ram_buffer(8956) := X"00000000";
		ram_buffer(8957) := X"00000000";
		ram_buffer(8958) := X"00000000";
		ram_buffer(8959) := X"00000000";
		ram_buffer(8960) := X"00000000";
		ram_buffer(8961) := X"00000000";
		ram_buffer(8962) := X"00000000";
		ram_buffer(8963) := X"00000000";
		ram_buffer(8964) := X"00000000";
		ram_buffer(8965) := X"00000000";
		ram_buffer(8966) := X"00000000";
		ram_buffer(8967) := X"00000000";
		ram_buffer(8968) := X"00000000";
		ram_buffer(8969) := X"00000000";
		ram_buffer(8970) := X"00000000";
		ram_buffer(8971) := X"00000000";
		ram_buffer(8972) := X"00000000";
		ram_buffer(8973) := X"00000000";
		ram_buffer(8974) := X"00000000";
		ram_buffer(8975) := X"00000000";
		ram_buffer(8976) := X"00000000";
		ram_buffer(8977) := X"00000000";
		ram_buffer(8978) := X"00000000";
		ram_buffer(8979) := X"00000000";
		ram_buffer(8980) := X"00000000";
		ram_buffer(8981) := X"00000000";
		ram_buffer(8982) := X"00000000";
		ram_buffer(8983) := X"00000000";
		ram_buffer(8984) := X"00000000";
		ram_buffer(8985) := X"00000000";
		ram_buffer(8986) := X"00000000";
		ram_buffer(8987) := X"00000000";
		ram_buffer(8988) := X"00000000";
		ram_buffer(8989) := X"00000000";
		ram_buffer(8990) := X"00000000";
		ram_buffer(8991) := X"00000000";
		ram_buffer(8992) := X"00000000";
		ram_buffer(8993) := X"00000000";
		ram_buffer(8994) := X"00000000";
		ram_buffer(8995) := X"00000000";
		ram_buffer(8996) := X"00000000";
		ram_buffer(8997) := X"00000000";
		ram_buffer(8998) := X"00000000";
		ram_buffer(8999) := X"00000000";
		ram_buffer(9000) := X"00000000";
		ram_buffer(9001) := X"00000000";
		ram_buffer(9002) := X"00000000";
		ram_buffer(9003) := X"00000000";
		ram_buffer(9004) := X"00000000";
		ram_buffer(9005) := X"00000000";
		ram_buffer(9006) := X"00000000";
		ram_buffer(9007) := X"00000000";
		ram_buffer(9008) := X"00000000";
		ram_buffer(9009) := X"00000000";
		ram_buffer(9010) := X"00000000";
		ram_buffer(9011) := X"00000000";
		ram_buffer(9012) := X"00000000";
		ram_buffer(9013) := X"00000000";
		ram_buffer(9014) := X"00000000";
		ram_buffer(9015) := X"00000000";
		ram_buffer(9016) := X"00000000";
		ram_buffer(9017) := X"00000000";
		ram_buffer(9018) := X"00000000";
		ram_buffer(9019) := X"00000000";
		ram_buffer(9020) := X"00000000";
		ram_buffer(9021) := X"00000000";
		ram_buffer(9022) := X"00000000";
		ram_buffer(9023) := X"00000000";
		ram_buffer(9024) := X"00000000";
		ram_buffer(9025) := X"00000000";
		ram_buffer(9026) := X"00000000";
		ram_buffer(9027) := X"00000000";
		ram_buffer(9028) := X"00000000";
		ram_buffer(9029) := X"00000000";
		ram_buffer(9030) := X"00000000";
		ram_buffer(9031) := X"00000000";
		ram_buffer(9032) := X"00000000";
		ram_buffer(9033) := X"00000000";
		ram_buffer(9034) := X"00000000";
		ram_buffer(9035) := X"00000000";
		ram_buffer(9036) := X"00000000";
		ram_buffer(9037) := X"00000000";
		ram_buffer(9038) := X"00000000";
		ram_buffer(9039) := X"00000000";
		ram_buffer(9040) := X"00000000";
		ram_buffer(9041) := X"00000000";
		ram_buffer(9042) := X"00000000";
		ram_buffer(9043) := X"00000000";
		ram_buffer(9044) := X"00000000";
		ram_buffer(9045) := X"00000000";
		ram_buffer(9046) := X"00000000";
		ram_buffer(9047) := X"00000000";
		ram_buffer(9048) := X"00000000";
		ram_buffer(9049) := X"00000000";
		ram_buffer(9050) := X"00000000";
		ram_buffer(9051) := X"00000000";
		ram_buffer(9052) := X"00000000";
		ram_buffer(9053) := X"00000000";
		ram_buffer(9054) := X"00000000";
		ram_buffer(9055) := X"00000000";
		ram_buffer(9056) := X"00000000";
		ram_buffer(9057) := X"00000000";
		ram_buffer(9058) := X"00000000";
		ram_buffer(9059) := X"00000000";
		ram_buffer(9060) := X"00000000";
		ram_buffer(9061) := X"00000000";
		ram_buffer(9062) := X"00000000";
		ram_buffer(9063) := X"00000000";
		ram_buffer(9064) := X"00000000";
		ram_buffer(9065) := X"00000000";
		ram_buffer(9066) := X"00000000";
		ram_buffer(9067) := X"00000000";
		ram_buffer(9068) := X"00000000";
		ram_buffer(9069) := X"00000000";
		ram_buffer(9070) := X"00000000";
		ram_buffer(9071) := X"00000000";
		ram_buffer(9072) := X"00000000";
		ram_buffer(9073) := X"00000000";
		ram_buffer(9074) := X"00000000";
		ram_buffer(9075) := X"00000000";
		ram_buffer(9076) := X"00000000";
		ram_buffer(9077) := X"00000000";
		ram_buffer(9078) := X"00000000";
		ram_buffer(9079) := X"00000000";
		ram_buffer(9080) := X"00000000";
		ram_buffer(9081) := X"00000000";
		ram_buffer(9082) := X"00000000";
		ram_buffer(9083) := X"00000000";
		ram_buffer(9084) := X"00000000";
		ram_buffer(9085) := X"00000000";
		ram_buffer(9086) := X"00000000";
		ram_buffer(9087) := X"00000000";
		ram_buffer(9088) := X"00000000";
		ram_buffer(9089) := X"00000000";
		ram_buffer(9090) := X"00000000";
		ram_buffer(9091) := X"00000000";
		ram_buffer(9092) := X"00000000";
		ram_buffer(9093) := X"00000000";
		ram_buffer(9094) := X"00000000";
		ram_buffer(9095) := X"00000000";
		ram_buffer(9096) := X"00000000";
		ram_buffer(9097) := X"00000000";
		ram_buffer(9098) := X"00000000";
		ram_buffer(9099) := X"00000000";
		ram_buffer(9100) := X"00000000";
		ram_buffer(9101) := X"00000000";
		ram_buffer(9102) := X"00000000";
		ram_buffer(9103) := X"00000000";
		ram_buffer(9104) := X"00000000";
		ram_buffer(9105) := X"00000000";
		ram_buffer(9106) := X"00000000";
		ram_buffer(9107) := X"00000000";
		ram_buffer(9108) := X"00000000";
		ram_buffer(9109) := X"00000000";
		ram_buffer(9110) := X"00000000";
		ram_buffer(9111) := X"00000000";
		ram_buffer(9112) := X"00000000";
		ram_buffer(9113) := X"00000000";
		ram_buffer(9114) := X"00000000";
		ram_buffer(9115) := X"00000000";
		ram_buffer(9116) := X"00000000";
		ram_buffer(9117) := X"00000000";
		ram_buffer(9118) := X"00000000";
		ram_buffer(9119) := X"00000000";
		ram_buffer(9120) := X"00000000";
		ram_buffer(9121) := X"00000000";
		ram_buffer(9122) := X"00000000";
		ram_buffer(9123) := X"00000000";
		ram_buffer(9124) := X"00000000";
		ram_buffer(9125) := X"00000000";
		ram_buffer(9126) := X"00000000";
		ram_buffer(9127) := X"00000000";
		ram_buffer(9128) := X"00000000";
		ram_buffer(9129) := X"00000000";
		ram_buffer(9130) := X"00000000";
		ram_buffer(9131) := X"00000000";
		ram_buffer(9132) := X"00000000";
		ram_buffer(9133) := X"00000000";
		ram_buffer(9134) := X"00000000";
		ram_buffer(9135) := X"00000000";
		ram_buffer(9136) := X"00000000";
		ram_buffer(9137) := X"00000000";
		ram_buffer(9138) := X"00000000";
		ram_buffer(9139) := X"00000000";
		ram_buffer(9140) := X"00000000";
		ram_buffer(9141) := X"00000000";
		ram_buffer(9142) := X"00000000";
		ram_buffer(9143) := X"00000000";
		ram_buffer(9144) := X"00000000";
		ram_buffer(9145) := X"00000000";
		ram_buffer(9146) := X"00000000";
		ram_buffer(9147) := X"00000000";
		ram_buffer(9148) := X"00000000";
		ram_buffer(9149) := X"00000000";
		ram_buffer(9150) := X"00000000";
		ram_buffer(9151) := X"00000000";
		ram_buffer(9152) := X"00000000";
		ram_buffer(9153) := X"00000000";
		ram_buffer(9154) := X"00000000";
		ram_buffer(9155) := X"00000000";
		ram_buffer(9156) := X"00000000";
		ram_buffer(9157) := X"00000000";
		ram_buffer(9158) := X"00000000";
		ram_buffer(9159) := X"00000000";
		ram_buffer(9160) := X"00000000";
		ram_buffer(9161) := X"00000000";
		ram_buffer(9162) := X"00000000";
		ram_buffer(9163) := X"00000000";
		ram_buffer(9164) := X"00000000";
		ram_buffer(9165) := X"00000000";
		ram_buffer(9166) := X"00000000";
		ram_buffer(9167) := X"00000000";
		ram_buffer(9168) := X"00000000";
		ram_buffer(9169) := X"00000000";
		ram_buffer(9170) := X"00000000";
		ram_buffer(9171) := X"00000000";
		ram_buffer(9172) := X"00000000";
		ram_buffer(9173) := X"00000000";
		ram_buffer(9174) := X"00000000";
		ram_buffer(9175) := X"00000000";
		ram_buffer(9176) := X"00000000";
		ram_buffer(9177) := X"00000000";
		ram_buffer(9178) := X"00000000";
		ram_buffer(9179) := X"00000000";
		ram_buffer(9180) := X"00000000";
		ram_buffer(9181) := X"00000000";
		ram_buffer(9182) := X"00000000";
		ram_buffer(9183) := X"00000000";
		ram_buffer(9184) := X"00000000";
		ram_buffer(9185) := X"00000000";
		ram_buffer(9186) := X"00000000";
		ram_buffer(9187) := X"00000000";
		ram_buffer(9188) := X"00000000";
		ram_buffer(9189) := X"00000000";
		ram_buffer(9190) := X"00000000";
		ram_buffer(9191) := X"00000000";
		ram_buffer(9192) := X"00000000";
		ram_buffer(9193) := X"00000000";
		ram_buffer(9194) := X"00000000";
		ram_buffer(9195) := X"00000000";
		ram_buffer(9196) := X"00000000";
		ram_buffer(9197) := X"00000000";
		ram_buffer(9198) := X"00000000";
		ram_buffer(9199) := X"00000000";
		ram_buffer(9200) := X"00000000";
		ram_buffer(9201) := X"00000000";
		ram_buffer(9202) := X"00000000";
		ram_buffer(9203) := X"00000000";
		ram_buffer(9204) := X"00000000";
		ram_buffer(9205) := X"00000000";
		ram_buffer(9206) := X"00000000";
		ram_buffer(9207) := X"00000000";
		ram_buffer(9208) := X"00000000";
		ram_buffer(9209) := X"00000000";
		ram_buffer(9210) := X"00000000";
		ram_buffer(9211) := X"00000000";
		ram_buffer(9212) := X"00000000";
		ram_buffer(9213) := X"00000000";
		ram_buffer(9214) := X"00000000";
		ram_buffer(9215) := X"00000000";
		ram_buffer(9216) := X"00000000";
		ram_buffer(9217) := X"00000000";
		ram_buffer(9218) := X"00000000";
		ram_buffer(9219) := X"00000000";
		ram_buffer(9220) := X"00000000";
		ram_buffer(9221) := X"00000000";
		ram_buffer(9222) := X"00000000";
		ram_buffer(9223) := X"00000000";
		ram_buffer(9224) := X"00000000";
		ram_buffer(9225) := X"00000000";
		ram_buffer(9226) := X"00000000";
		ram_buffer(9227) := X"00000000";
		ram_buffer(9228) := X"00000000";
		ram_buffer(9229) := X"00000000";
		ram_buffer(9230) := X"00000000";
		ram_buffer(9231) := X"00000000";
		ram_buffer(9232) := X"00000000";
		ram_buffer(9233) := X"00000000";
		ram_buffer(9234) := X"00000000";
		ram_buffer(9235) := X"00000000";
		ram_buffer(9236) := X"00000000";
		ram_buffer(9237) := X"00000000";
		ram_buffer(9238) := X"00000000";
		ram_buffer(9239) := X"00000000";
		ram_buffer(9240) := X"00000000";
		ram_buffer(9241) := X"00000000";
		ram_buffer(9242) := X"00000000";
		ram_buffer(9243) := X"00000000";
		ram_buffer(9244) := X"00000000";
		ram_buffer(9245) := X"00000000";
		ram_buffer(9246) := X"00000000";
		ram_buffer(9247) := X"00000000";
		ram_buffer(9248) := X"00000000";
		ram_buffer(9249) := X"00000000";
		ram_buffer(9250) := X"00000000";
		ram_buffer(9251) := X"00000000";
		ram_buffer(9252) := X"00000000";
		ram_buffer(9253) := X"00000000";
		ram_buffer(9254) := X"00000000";
		ram_buffer(9255) := X"00000000";
		ram_buffer(9256) := X"00000000";
		ram_buffer(9257) := X"00000000";
		ram_buffer(9258) := X"00000000";
		ram_buffer(9259) := X"00000000";
		ram_buffer(9260) := X"00000000";
		ram_buffer(9261) := X"00000000";
		ram_buffer(9262) := X"00000000";
		ram_buffer(9263) := X"00000000";
		ram_buffer(9264) := X"00000000";
		ram_buffer(9265) := X"00000000";
		ram_buffer(9266) := X"00000000";
		ram_buffer(9267) := X"00000000";
		ram_buffer(9268) := X"00000000";
		ram_buffer(9269) := X"00000000";
		ram_buffer(9270) := X"00000000";
		ram_buffer(9271) := X"00000000";
		ram_buffer(9272) := X"00000000";
		ram_buffer(9273) := X"00000000";
		ram_buffer(9274) := X"00000000";
		ram_buffer(9275) := X"00000000";
		ram_buffer(9276) := X"00000000";
		ram_buffer(9277) := X"00000000";
		ram_buffer(9278) := X"00000000";
		ram_buffer(9279) := X"00000000";
		ram_buffer(9280) := X"00000000";
		ram_buffer(9281) := X"00000000";
		ram_buffer(9282) := X"00000000";
		ram_buffer(9283) := X"00000000";
		ram_buffer(9284) := X"00000000";
		ram_buffer(9285) := X"00000000";
		ram_buffer(9286) := X"00000000";
		ram_buffer(9287) := X"00000000";
		ram_buffer(9288) := X"00000000";
		ram_buffer(9289) := X"00000000";
		ram_buffer(9290) := X"00000000";
		ram_buffer(9291) := X"00000000";
		ram_buffer(9292) := X"00000000";
		ram_buffer(9293) := X"00000000";
		ram_buffer(9294) := X"00000000";
		ram_buffer(9295) := X"00000000";
		ram_buffer(9296) := X"00000000";
		ram_buffer(9297) := X"00000000";
		ram_buffer(9298) := X"00000000";
		ram_buffer(9299) := X"00000000";
		ram_buffer(9300) := X"00000000";
		ram_buffer(9301) := X"00000000";
		ram_buffer(9302) := X"00000000";
		ram_buffer(9303) := X"00000000";
		ram_buffer(9304) := X"00000000";
		ram_buffer(9305) := X"00000000";
		ram_buffer(9306) := X"00000000";
		ram_buffer(9307) := X"00000000";
		ram_buffer(9308) := X"00000000";
		ram_buffer(9309) := X"00000000";
		ram_buffer(9310) := X"00000000";
		ram_buffer(9311) := X"00000000";
		ram_buffer(9312) := X"00000000";
		ram_buffer(9313) := X"00000000";
		ram_buffer(9314) := X"00000000";
		ram_buffer(9315) := X"00000000";
		ram_buffer(9316) := X"00000000";
		ram_buffer(9317) := X"00000000";
		ram_buffer(9318) := X"00000000";
		ram_buffer(9319) := X"00000000";
		ram_buffer(9320) := X"00000000";
		ram_buffer(9321) := X"00000000";
		ram_buffer(9322) := X"00000000";
		ram_buffer(9323) := X"00000000";
		ram_buffer(9324) := X"00000000";
		ram_buffer(9325) := X"00000000";
		ram_buffer(9326) := X"00000000";
		ram_buffer(9327) := X"00000000";
		ram_buffer(9328) := X"00000000";
		ram_buffer(9329) := X"00000000";
		ram_buffer(9330) := X"00000000";
		ram_buffer(9331) := X"00000000";
		ram_buffer(9332) := X"00000000";
		ram_buffer(9333) := X"00000000";
		ram_buffer(9334) := X"00000000";
		ram_buffer(9335) := X"00000000";
		ram_buffer(9336) := X"00000000";
		ram_buffer(9337) := X"00000000";
		ram_buffer(9338) := X"00000000";
		ram_buffer(9339) := X"00000000";
		ram_buffer(9340) := X"00000000";
		ram_buffer(9341) := X"00000000";
		ram_buffer(9342) := X"00000000";
		ram_buffer(9343) := X"00000000";
		ram_buffer(9344) := X"00000000";
		ram_buffer(9345) := X"00000000";
		ram_buffer(9346) := X"00000000";
		ram_buffer(9347) := X"00000000";
		ram_buffer(9348) := X"00000000";
		ram_buffer(9349) := X"00000000";
		ram_buffer(9350) := X"00000000";
		ram_buffer(9351) := X"00000000";
		ram_buffer(9352) := X"00000000";
		ram_buffer(9353) := X"00000000";
		ram_buffer(9354) := X"00000000";
		ram_buffer(9355) := X"00000000";
		ram_buffer(9356) := X"00000000";
		ram_buffer(9357) := X"00000000";
		ram_buffer(9358) := X"00000000";
		ram_buffer(9359) := X"00000000";
		ram_buffer(9360) := X"00000000";
		ram_buffer(9361) := X"00000000";
		ram_buffer(9362) := X"00000000";
		ram_buffer(9363) := X"00000000";
		ram_buffer(9364) := X"00000000";
		ram_buffer(9365) := X"00000000";
		ram_buffer(9366) := X"00000000";
		ram_buffer(9367) := X"00000000";
		ram_buffer(9368) := X"00000000";
		ram_buffer(9369) := X"00000000";
		ram_buffer(9370) := X"00000000";
		ram_buffer(9371) := X"00000000";
		ram_buffer(9372) := X"00000000";
		ram_buffer(9373) := X"00000000";
		ram_buffer(9374) := X"00000000";
		ram_buffer(9375) := X"00000000";
		ram_buffer(9376) := X"00000000";
		ram_buffer(9377) := X"00000000";
		ram_buffer(9378) := X"00000000";
		ram_buffer(9379) := X"00000000";
		ram_buffer(9380) := X"00000000";
		ram_buffer(9381) := X"00000000";
		ram_buffer(9382) := X"00000000";
		ram_buffer(9383) := X"00000000";
		ram_buffer(9384) := X"00000000";
		ram_buffer(9385) := X"00000000";
		ram_buffer(9386) := X"00000000";
		ram_buffer(9387) := X"00000000";
		ram_buffer(9388) := X"00000000";
		ram_buffer(9389) := X"00000000";
		ram_buffer(9390) := X"00000000";
		ram_buffer(9391) := X"00000000";
		ram_buffer(9392) := X"00000000";
		ram_buffer(9393) := X"00000000";
		ram_buffer(9394) := X"00000000";
		ram_buffer(9395) := X"00000000";
		ram_buffer(9396) := X"00000000";
		ram_buffer(9397) := X"00000000";
		ram_buffer(9398) := X"00000000";
		ram_buffer(9399) := X"00000000";
		ram_buffer(9400) := X"00000000";
		ram_buffer(9401) := X"00000000";
		ram_buffer(9402) := X"00000000";
		ram_buffer(9403) := X"00000000";
		ram_buffer(9404) := X"00000000";
		ram_buffer(9405) := X"00000000";
		ram_buffer(9406) := X"00000000";
		ram_buffer(9407) := X"00000000";
		ram_buffer(9408) := X"00000000";
		ram_buffer(9409) := X"00000000";
		ram_buffer(9410) := X"00000000";
		ram_buffer(9411) := X"00000000";
		ram_buffer(9412) := X"00000000";
		ram_buffer(9413) := X"00000000";
		ram_buffer(9414) := X"00000000";
		ram_buffer(9415) := X"00000000";
		ram_buffer(9416) := X"00000000";
		ram_buffer(9417) := X"00000000";
		ram_buffer(9418) := X"00000000";
		ram_buffer(9419) := X"00000000";
		ram_buffer(9420) := X"00000000";
		ram_buffer(9421) := X"00000000";
		ram_buffer(9422) := X"00000000";
		ram_buffer(9423) := X"00000000";
		ram_buffer(9424) := X"00000000";
		ram_buffer(9425) := X"00000000";
		ram_buffer(9426) := X"00000000";
		ram_buffer(9427) := X"00000000";
		ram_buffer(9428) := X"00000000";
		ram_buffer(9429) := X"00000000";
		ram_buffer(9430) := X"00000000";
		ram_buffer(9431) := X"00000000";
		ram_buffer(9432) := X"00000000";
		ram_buffer(9433) := X"00000000";
		ram_buffer(9434) := X"00000000";
		ram_buffer(9435) := X"00000000";
		ram_buffer(9436) := X"00000000";
		ram_buffer(9437) := X"00000000";
		ram_buffer(9438) := X"00000000";
		ram_buffer(9439) := X"00000000";
		ram_buffer(9440) := X"00000000";
		ram_buffer(9441) := X"00000000";
		ram_buffer(9442) := X"00000000";
		ram_buffer(9443) := X"00000000";
		ram_buffer(9444) := X"00000000";
		ram_buffer(9445) := X"00000000";
		ram_buffer(9446) := X"00000000";
		ram_buffer(9447) := X"00000000";
		ram_buffer(9448) := X"00000000";
		ram_buffer(9449) := X"00000000";
		ram_buffer(9450) := X"00000000";
		ram_buffer(9451) := X"00000000";
		ram_buffer(9452) := X"00000000";
		ram_buffer(9453) := X"00000000";
		ram_buffer(9454) := X"00000000";
		ram_buffer(9455) := X"00000000";
		ram_buffer(9456) := X"00000000";
		ram_buffer(9457) := X"00000000";
		ram_buffer(9458) := X"00000000";
		ram_buffer(9459) := X"00000000";
		ram_buffer(9460) := X"00000000";
		ram_buffer(9461) := X"00000000";
		ram_buffer(9462) := X"00000000";
		ram_buffer(9463) := X"00000000";
		ram_buffer(9464) := X"00000000";
		ram_buffer(9465) := X"00000000";
		ram_buffer(9466) := X"00000000";
		ram_buffer(9467) := X"00000000";
		ram_buffer(9468) := X"00000000";
		ram_buffer(9469) := X"00000000";
		ram_buffer(9470) := X"00000000";
		ram_buffer(9471) := X"00000000";
		ram_buffer(9472) := X"00000000";
		ram_buffer(9473) := X"00000000";
		ram_buffer(9474) := X"00000000";
		ram_buffer(9475) := X"00000000";
		ram_buffer(9476) := X"00000000";
		ram_buffer(9477) := X"00000000";
		ram_buffer(9478) := X"00000000";
		ram_buffer(9479) := X"00000000";
		ram_buffer(9480) := X"00000000";
		ram_buffer(9481) := X"00000000";
		ram_buffer(9482) := X"00000000";
		ram_buffer(9483) := X"00000000";
		ram_buffer(9484) := X"00000000";
		ram_buffer(9485) := X"00000000";
		ram_buffer(9486) := X"00000000";
		ram_buffer(9487) := X"00000000";
		ram_buffer(9488) := X"00000000";
		ram_buffer(9489) := X"00000000";
		ram_buffer(9490) := X"00000000";
		ram_buffer(9491) := X"00000000";
		ram_buffer(9492) := X"00000000";
		ram_buffer(9493) := X"00000000";
		ram_buffer(9494) := X"00000000";
		ram_buffer(9495) := X"00000000";
		ram_buffer(9496) := X"00000000";
		ram_buffer(9497) := X"00000000";
		ram_buffer(9498) := X"00000000";
		ram_buffer(9499) := X"00000000";
		ram_buffer(9500) := X"00000000";
		ram_buffer(9501) := X"00000000";
		ram_buffer(9502) := X"00000000";
		ram_buffer(9503) := X"00000000";
		ram_buffer(9504) := X"00000000";
		ram_buffer(9505) := X"00000000";
		ram_buffer(9506) := X"00000000";
		ram_buffer(9507) := X"00000000";
		ram_buffer(9508) := X"00000000";
		ram_buffer(9509) := X"00000000";
		ram_buffer(9510) := X"00000000";
		ram_buffer(9511) := X"00000000";
		ram_buffer(9512) := X"00000000";
		ram_buffer(9513) := X"00000000";
		ram_buffer(9514) := X"00000000";
		ram_buffer(9515) := X"00000000";
		ram_buffer(9516) := X"00000000";
		ram_buffer(9517) := X"00000000";
		ram_buffer(9518) := X"00000000";
		ram_buffer(9519) := X"00000000";
		ram_buffer(9520) := X"00000000";
		ram_buffer(9521) := X"00000000";
		ram_buffer(9522) := X"00000000";
		ram_buffer(9523) := X"00000000";
		ram_buffer(9524) := X"00000000";
		ram_buffer(9525) := X"00000000";
		ram_buffer(9526) := X"00000000";
		ram_buffer(9527) := X"00000000";
		ram_buffer(9528) := X"00000000";
		ram_buffer(9529) := X"00000000";
		ram_buffer(9530) := X"00000000";
		ram_buffer(9531) := X"00000000";
		ram_buffer(9532) := X"00000000";
		ram_buffer(9533) := X"00000000";
		ram_buffer(9534) := X"00000000";
		ram_buffer(9535) := X"00000000";
		ram_buffer(9536) := X"00000000";
		ram_buffer(9537) := X"00000000";
		ram_buffer(9538) := X"00000000";
		ram_buffer(9539) := X"00000000";
		ram_buffer(9540) := X"00000000";
		ram_buffer(9541) := X"00000000";
		ram_buffer(9542) := X"00000000";
		ram_buffer(9543) := X"00000000";
		ram_buffer(9544) := X"00000000";
		ram_buffer(9545) := X"00000000";
		ram_buffer(9546) := X"00000000";
		ram_buffer(9547) := X"00000000";
		ram_buffer(9548) := X"00000000";
		ram_buffer(9549) := X"00000000";
		ram_buffer(9550) := X"00000000";
		ram_buffer(9551) := X"00000000";
		ram_buffer(9552) := X"00000000";
		ram_buffer(9553) := X"00000000";
		ram_buffer(9554) := X"00000000";
		ram_buffer(9555) := X"00000000";
		ram_buffer(9556) := X"00000000";
		ram_buffer(9557) := X"00000000";
		ram_buffer(9558) := X"00000000";
		ram_buffer(9559) := X"00000000";
		ram_buffer(9560) := X"00000000";
		ram_buffer(9561) := X"00000000";
		ram_buffer(9562) := X"00000000";
		ram_buffer(9563) := X"00000000";
		ram_buffer(9564) := X"00000000";
		ram_buffer(9565) := X"00000000";
		ram_buffer(9566) := X"00000000";
		ram_buffer(9567) := X"00000000";
		ram_buffer(9568) := X"00000000";
		ram_buffer(9569) := X"00000000";
		ram_buffer(9570) := X"00000000";
		ram_buffer(9571) := X"00000000";
		ram_buffer(9572) := X"00000000";
		ram_buffer(9573) := X"00000000";
		ram_buffer(9574) := X"00000000";
		ram_buffer(9575) := X"00000000";
		ram_buffer(9576) := X"00000000";
		ram_buffer(9577) := X"00000000";
		ram_buffer(9578) := X"00000000";
		ram_buffer(9579) := X"00000000";
		ram_buffer(9580) := X"00000000";
		ram_buffer(9581) := X"00000000";
		ram_buffer(9582) := X"00000000";
		ram_buffer(9583) := X"00000000";
		ram_buffer(9584) := X"00000000";
		ram_buffer(9585) := X"00000000";
		ram_buffer(9586) := X"00000000";
		ram_buffer(9587) := X"00000000";
		ram_buffer(9588) := X"00000000";
		ram_buffer(9589) := X"00000000";
		ram_buffer(9590) := X"00000000";
		ram_buffer(9591) := X"00000000";
		ram_buffer(9592) := X"00000000";
		ram_buffer(9593) := X"00000000";
		ram_buffer(9594) := X"00000000";
		ram_buffer(9595) := X"00000000";
		ram_buffer(9596) := X"00000000";
		ram_buffer(9597) := X"00000000";
		ram_buffer(9598) := X"00000000";
		ram_buffer(9599) := X"00000000";
		ram_buffer(9600) := X"00000000";
		ram_buffer(9601) := X"00000000";
		ram_buffer(9602) := X"00000000";
		ram_buffer(9603) := X"00000000";
		ram_buffer(9604) := X"00000000";
		ram_buffer(9605) := X"00000000";
		ram_buffer(9606) := X"00000000";
		ram_buffer(9607) := X"00000000";
		ram_buffer(9608) := X"00000000";
		ram_buffer(9609) := X"00000000";
		ram_buffer(9610) := X"00000000";
		ram_buffer(9611) := X"00000000";
		ram_buffer(9612) := X"00000000";
		ram_buffer(9613) := X"00000000";
		ram_buffer(9614) := X"00000000";
		ram_buffer(9615) := X"00000000";
		ram_buffer(9616) := X"00000000";
		ram_buffer(9617) := X"00000000";
		ram_buffer(9618) := X"00000000";
		ram_buffer(9619) := X"00000000";
		ram_buffer(9620) := X"00000000";
		ram_buffer(9621) := X"00000000";
		ram_buffer(9622) := X"00000000";
		ram_buffer(9623) := X"00000000";
		ram_buffer(9624) := X"00000000";
		ram_buffer(9625) := X"00000000";
		ram_buffer(9626) := X"00000000";
		ram_buffer(9627) := X"00000000";
		ram_buffer(9628) := X"00000000";
		ram_buffer(9629) := X"00000000";
		ram_buffer(9630) := X"00000000";
		ram_buffer(9631) := X"00000000";
		ram_buffer(9632) := X"00000000";
		ram_buffer(9633) := X"00000000";
		ram_buffer(9634) := X"00000000";
		ram_buffer(9635) := X"00000000";
		ram_buffer(9636) := X"00000000";
		ram_buffer(9637) := X"00000000";
		ram_buffer(9638) := X"00000000";
		ram_buffer(9639) := X"00000000";
		ram_buffer(9640) := X"00000000";
		ram_buffer(9641) := X"00000000";
		ram_buffer(9642) := X"00000000";
		ram_buffer(9643) := X"00000000";
		ram_buffer(9644) := X"00000000";
		ram_buffer(9645) := X"00000000";
		ram_buffer(9646) := X"00000000";
		ram_buffer(9647) := X"00000000";
		ram_buffer(9648) := X"00000000";
		ram_buffer(9649) := X"00000000";
		ram_buffer(9650) := X"00000000";
		ram_buffer(9651) := X"00000000";
		ram_buffer(9652) := X"00000000";
		ram_buffer(9653) := X"00000000";
		ram_buffer(9654) := X"00000000";
		ram_buffer(9655) := X"00000000";
		ram_buffer(9656) := X"00000000";
		ram_buffer(9657) := X"00000000";
		ram_buffer(9658) := X"00000000";
		ram_buffer(9659) := X"00000000";
		ram_buffer(9660) := X"00000000";
		ram_buffer(9661) := X"00000000";
		ram_buffer(9662) := X"00000000";
		ram_buffer(9663) := X"00000000";
		ram_buffer(9664) := X"00000000";
		ram_buffer(9665) := X"00000000";
		ram_buffer(9666) := X"00000000";
		ram_buffer(9667) := X"00000000";
		ram_buffer(9668) := X"00000000";
		ram_buffer(9669) := X"00000000";
		ram_buffer(9670) := X"00000000";
		ram_buffer(9671) := X"00000000";
		ram_buffer(9672) := X"00000000";
		ram_buffer(9673) := X"00000000";
		ram_buffer(9674) := X"00000000";
		ram_buffer(9675) := X"00000000";
		ram_buffer(9676) := X"00000000";
		ram_buffer(9677) := X"00000000";
		ram_buffer(9678) := X"00000000";
		ram_buffer(9679) := X"00000000";
		ram_buffer(9680) := X"00000000";
		ram_buffer(9681) := X"00000000";
		ram_buffer(9682) := X"00000000";
		ram_buffer(9683) := X"00000000";
		ram_buffer(9684) := X"00000000";
		ram_buffer(9685) := X"00000000";
		ram_buffer(9686) := X"00000000";
		ram_buffer(9687) := X"00000000";
		ram_buffer(9688) := X"00000000";
		ram_buffer(9689) := X"00000000";
		ram_buffer(9690) := X"00000000";
		ram_buffer(9691) := X"00000000";
		ram_buffer(9692) := X"00000000";
		ram_buffer(9693) := X"00000000";
		ram_buffer(9694) := X"00000000";
		ram_buffer(9695) := X"00000000";
		ram_buffer(9696) := X"00000000";
		ram_buffer(9697) := X"00000000";
		ram_buffer(9698) := X"00000000";
		ram_buffer(9699) := X"00000000";
		ram_buffer(9700) := X"00000000";
		ram_buffer(9701) := X"00000000";
		ram_buffer(9702) := X"00000000";
		ram_buffer(9703) := X"00000000";
		ram_buffer(9704) := X"00000000";
		ram_buffer(9705) := X"00000000";
		ram_buffer(9706) := X"00000000";
		ram_buffer(9707) := X"00000000";
		ram_buffer(9708) := X"00000000";
		ram_buffer(9709) := X"00000000";
		ram_buffer(9710) := X"00000000";
		ram_buffer(9711) := X"00000000";
		ram_buffer(9712) := X"00000000";
		ram_buffer(9713) := X"00000000";
		ram_buffer(9714) := X"00000000";
		ram_buffer(9715) := X"00000000";
		ram_buffer(9716) := X"00000000";
		ram_buffer(9717) := X"00000000";
		ram_buffer(9718) := X"00000000";
		ram_buffer(9719) := X"00000000";
		ram_buffer(9720) := X"00000000";
		ram_buffer(9721) := X"00000000";
		ram_buffer(9722) := X"00000000";
		ram_buffer(9723) := X"00000000";
		ram_buffer(9724) := X"00000000";
		ram_buffer(9725) := X"00000000";
		ram_buffer(9726) := X"00000000";
		ram_buffer(9727) := X"00000000";
		ram_buffer(9728) := X"00000000";
		ram_buffer(9729) := X"00000000";
		ram_buffer(9730) := X"00000000";
		ram_buffer(9731) := X"00000000";
		ram_buffer(9732) := X"00000000";
		ram_buffer(9733) := X"00000000";
		ram_buffer(9734) := X"00000000";
		ram_buffer(9735) := X"00000000";
		ram_buffer(9736) := X"00000000";
		ram_buffer(9737) := X"00000000";
		ram_buffer(9738) := X"00000000";
		ram_buffer(9739) := X"00000000";
		ram_buffer(9740) := X"00000000";
		ram_buffer(9741) := X"00000000";
		ram_buffer(9742) := X"00000000";
		ram_buffer(9743) := X"00000000";
		ram_buffer(9744) := X"00000000";
		ram_buffer(9745) := X"00000000";
		ram_buffer(9746) := X"00000000";
		ram_buffer(9747) := X"00000000";
		ram_buffer(9748) := X"00000000";
		ram_buffer(9749) := X"00000000";
		ram_buffer(9750) := X"00000000";
		ram_buffer(9751) := X"00000000";
		ram_buffer(9752) := X"00000000";
		ram_buffer(9753) := X"00000000";
		ram_buffer(9754) := X"00000000";
		ram_buffer(9755) := X"00000000";
		ram_buffer(9756) := X"00000000";
		ram_buffer(9757) := X"00000000";
		ram_buffer(9758) := X"00000000";
		ram_buffer(9759) := X"00000000";
		ram_buffer(9760) := X"00000000";
		ram_buffer(9761) := X"00000000";
		ram_buffer(9762) := X"00000000";
		ram_buffer(9763) := X"00000000";
		ram_buffer(9764) := X"00000000";
		ram_buffer(9765) := X"00000000";
		ram_buffer(9766) := X"00000000";
		ram_buffer(9767) := X"00000000";
		ram_buffer(9768) := X"00000000";
		ram_buffer(9769) := X"00000000";
		ram_buffer(9770) := X"00000000";
		ram_buffer(9771) := X"00000000";
		ram_buffer(9772) := X"00000000";
		ram_buffer(9773) := X"00000000";
		ram_buffer(9774) := X"00000000";
		ram_buffer(9775) := X"00000000";
		ram_buffer(9776) := X"00000000";
		ram_buffer(9777) := X"00000000";
		ram_buffer(9778) := X"00000000";
		ram_buffer(9779) := X"00000000";
		ram_buffer(9780) := X"00000000";
		ram_buffer(9781) := X"00000000";
		ram_buffer(9782) := X"00000000";
		ram_buffer(9783) := X"00000000";
		ram_buffer(9784) := X"00000000";
		ram_buffer(9785) := X"00000000";
		ram_buffer(9786) := X"00000000";
		ram_buffer(9787) := X"00000000";
		ram_buffer(9788) := X"00000000";
		ram_buffer(9789) := X"00000000";
		ram_buffer(9790) := X"00000000";
		ram_buffer(9791) := X"00000000";
		ram_buffer(9792) := X"00000000";
		ram_buffer(9793) := X"00000000";
		ram_buffer(9794) := X"00000000";
		ram_buffer(9795) := X"00000000";
		ram_buffer(9796) := X"00000000";
		ram_buffer(9797) := X"00000000";
		ram_buffer(9798) := X"00000000";
		ram_buffer(9799) := X"00000000";
		ram_buffer(9800) := X"00000000";
		ram_buffer(9801) := X"00000000";
		ram_buffer(9802) := X"00000000";
		ram_buffer(9803) := X"00000000";
		ram_buffer(9804) := X"00000000";
		ram_buffer(9805) := X"00000000";
		ram_buffer(9806) := X"00000000";
		ram_buffer(9807) := X"00000000";
		ram_buffer(9808) := X"00000000";
		ram_buffer(9809) := X"00000000";
		ram_buffer(9810) := X"00000000";
		ram_buffer(9811) := X"00000000";
		ram_buffer(9812) := X"00000000";
		ram_buffer(9813) := X"00000000";
		ram_buffer(9814) := X"00000000";
		ram_buffer(9815) := X"00000000";
		ram_buffer(9816) := X"00000000";
		ram_buffer(9817) := X"00000000";
		ram_buffer(9818) := X"00000000";
		ram_buffer(9819) := X"00000000";
		ram_buffer(9820) := X"00000000";
		ram_buffer(9821) := X"00000000";
		ram_buffer(9822) := X"00000000";
		ram_buffer(9823) := X"00000000";
		ram_buffer(9824) := X"00000000";
		ram_buffer(9825) := X"00000000";
		ram_buffer(9826) := X"00000000";
		ram_buffer(9827) := X"00000000";
		ram_buffer(9828) := X"00000000";
		ram_buffer(9829) := X"00000000";
		ram_buffer(9830) := X"00000000";
		ram_buffer(9831) := X"00000000";
		ram_buffer(9832) := X"00000000";
		ram_buffer(9833) := X"00000000";
		ram_buffer(9834) := X"00000000";
		ram_buffer(9835) := X"00000000";
		ram_buffer(9836) := X"00000000";
		ram_buffer(9837) := X"00000000";
		ram_buffer(9838) := X"00000000";
		ram_buffer(9839) := X"00000000";
		ram_buffer(9840) := X"00000000";
		ram_buffer(9841) := X"00000000";
		ram_buffer(9842) := X"00000000";
		ram_buffer(9843) := X"00000000";
		ram_buffer(9844) := X"00000000";
		ram_buffer(9845) := X"00000000";
		ram_buffer(9846) := X"00000000";
		ram_buffer(9847) := X"00000000";
		ram_buffer(9848) := X"00000000";
		ram_buffer(9849) := X"00000000";
		ram_buffer(9850) := X"00000000";
		ram_buffer(9851) := X"00000000";
		ram_buffer(9852) := X"00000000";
		ram_buffer(9853) := X"00000000";
		ram_buffer(9854) := X"00000000";
		ram_buffer(9855) := X"00000000";
		ram_buffer(9856) := X"00000000";
		ram_buffer(9857) := X"00000000";
		ram_buffer(9858) := X"00000000";
		ram_buffer(9859) := X"00000000";
		ram_buffer(9860) := X"00000000";
		ram_buffer(9861) := X"00000000";
		ram_buffer(9862) := X"00000000";
		ram_buffer(9863) := X"00000000";
		ram_buffer(9864) := X"00000000";
		ram_buffer(9865) := X"00000000";
		ram_buffer(9866) := X"00000000";
		ram_buffer(9867) := X"00000000";
		ram_buffer(9868) := X"00000000";
		ram_buffer(9869) := X"00000000";
		ram_buffer(9870) := X"00000000";
		ram_buffer(9871) := X"00000000";
		ram_buffer(9872) := X"00000000";
		ram_buffer(9873) := X"00000000";
		ram_buffer(9874) := X"00000000";
		ram_buffer(9875) := X"00000000";
		ram_buffer(9876) := X"00000000";
		ram_buffer(9877) := X"00000000";
		ram_buffer(9878) := X"00000000";
		ram_buffer(9879) := X"00000000";
		ram_buffer(9880) := X"00000000";
		ram_buffer(9881) := X"00000000";
		ram_buffer(9882) := X"00000000";
		ram_buffer(9883) := X"00000000";
		ram_buffer(9884) := X"00000000";
		ram_buffer(9885) := X"00000000";
		ram_buffer(9886) := X"00000000";
		ram_buffer(9887) := X"00000000";
		ram_buffer(9888) := X"00000000";
		ram_buffer(9889) := X"00000000";
		ram_buffer(9890) := X"00000000";
		ram_buffer(9891) := X"00000000";
		ram_buffer(9892) := X"00000000";
		ram_buffer(9893) := X"00000000";
		ram_buffer(9894) := X"00000000";
		ram_buffer(9895) := X"00000000";
		ram_buffer(9896) := X"00000000";
		ram_buffer(9897) := X"00000000";
		ram_buffer(9898) := X"00000000";
		ram_buffer(9899) := X"00000000";
		ram_buffer(9900) := X"00000000";
		ram_buffer(9901) := X"00000000";
		ram_buffer(9902) := X"00000000";
		ram_buffer(9903) := X"00000000";
		ram_buffer(9904) := X"00000000";
		ram_buffer(9905) := X"00000000";
		ram_buffer(9906) := X"00000000";
		ram_buffer(9907) := X"00000000";
		ram_buffer(9908) := X"00000000";
		ram_buffer(9909) := X"00000000";
		ram_buffer(9910) := X"00000000";
		ram_buffer(9911) := X"00000000";
		ram_buffer(9912) := X"00000000";
		ram_buffer(9913) := X"00000000";
		ram_buffer(9914) := X"00000000";
		ram_buffer(9915) := X"00000000";
		ram_buffer(9916) := X"00000000";
		ram_buffer(9917) := X"00000000";
		ram_buffer(9918) := X"00000000";
		ram_buffer(9919) := X"00000000";
		ram_buffer(9920) := X"00000000";
		ram_buffer(9921) := X"00000000";
		ram_buffer(9922) := X"00000000";
		ram_buffer(9923) := X"00000000";
		ram_buffer(9924) := X"00000000";
		ram_buffer(9925) := X"00000000";
		ram_buffer(9926) := X"00000000";
		ram_buffer(9927) := X"00000000";
		ram_buffer(9928) := X"00000000";
		ram_buffer(9929) := X"00000000";
		ram_buffer(9930) := X"00000000";
		ram_buffer(9931) := X"00000000";
		ram_buffer(9932) := X"00000000";
		ram_buffer(9933) := X"00000000";
		ram_buffer(9934) := X"00000000";
		ram_buffer(9935) := X"00000000";
		ram_buffer(9936) := X"00000000";
		ram_buffer(9937) := X"00000000";
		ram_buffer(9938) := X"00000000";
		ram_buffer(9939) := X"00000000";
		ram_buffer(9940) := X"00000000";
		ram_buffer(9941) := X"00000000";
		ram_buffer(9942) := X"00000000";
		ram_buffer(9943) := X"00000000";
		ram_buffer(9944) := X"00000000";
		ram_buffer(9945) := X"00000000";
		ram_buffer(9946) := X"00000000";
		ram_buffer(9947) := X"00000000";
		ram_buffer(9948) := X"00000000";
		ram_buffer(9949) := X"00000000";
		ram_buffer(9950) := X"00000000";
		ram_buffer(9951) := X"00000000";
		ram_buffer(9952) := X"00000000";
		ram_buffer(9953) := X"00000000";
		ram_buffer(9954) := X"00000000";
		ram_buffer(9955) := X"00000000";
		ram_buffer(9956) := X"00000000";
		ram_buffer(9957) := X"00000000";
		ram_buffer(9958) := X"00000000";
		ram_buffer(9959) := X"00000000";
		ram_buffer(9960) := X"00000000";
		ram_buffer(9961) := X"00000000";
		ram_buffer(9962) := X"00000000";
		ram_buffer(9963) := X"00000000";
		ram_buffer(9964) := X"00000000";
		ram_buffer(9965) := X"00000000";
		ram_buffer(9966) := X"00000000";
		ram_buffer(9967) := X"00000000";
		ram_buffer(9968) := X"00000000";
		ram_buffer(9969) := X"00000000";
		ram_buffer(9970) := X"00000000";
		ram_buffer(9971) := X"00000000";
		ram_buffer(9972) := X"00000000";
		ram_buffer(9973) := X"00000000";
		ram_buffer(9974) := X"00000000";
		ram_buffer(9975) := X"00000000";
		ram_buffer(9976) := X"00000000";
		ram_buffer(9977) := X"00000000";
		ram_buffer(9978) := X"00000000";
		ram_buffer(9979) := X"00000000";
		ram_buffer(9980) := X"00000000";
		ram_buffer(9981) := X"00000000";
		ram_buffer(9982) := X"00000000";
		ram_buffer(9983) := X"00000000";
		ram_buffer(9984) := X"00000000";
		ram_buffer(9985) := X"00000000";
		ram_buffer(9986) := X"00000000";
		ram_buffer(9987) := X"00000000";
		ram_buffer(9988) := X"00000000";
		ram_buffer(9989) := X"00000000";
		ram_buffer(9990) := X"00000000";
		ram_buffer(9991) := X"00000000";
		ram_buffer(9992) := X"00000000";
		ram_buffer(9993) := X"00000000";
		ram_buffer(9994) := X"00000000";
		ram_buffer(9995) := X"00000000";
		ram_buffer(9996) := X"00000000";
		ram_buffer(9997) := X"00000000";
		ram_buffer(9998) := X"00000000";
		ram_buffer(9999) := X"00000000";
		ram_buffer(10000) := X"00000000";
		ram_buffer(10001) := X"00000000";
		ram_buffer(10002) := X"00000000";
		ram_buffer(10003) := X"00000000";
		ram_buffer(10004) := X"00000000";
		ram_buffer(10005) := X"00000000";
		ram_buffer(10006) := X"00000000";
		ram_buffer(10007) := X"00000000";
		ram_buffer(10008) := X"00000000";
		ram_buffer(10009) := X"00000000";
		ram_buffer(10010) := X"00000000";
		ram_buffer(10011) := X"00000000";
		ram_buffer(10012) := X"00000000";
		ram_buffer(10013) := X"00000000";
		ram_buffer(10014) := X"00000000";
		ram_buffer(10015) := X"00000000";
		ram_buffer(10016) := X"00000000";
		ram_buffer(10017) := X"00000000";
		ram_buffer(10018) := X"00000000";
		ram_buffer(10019) := X"00000000";
		ram_buffer(10020) := X"00000000";
		ram_buffer(10021) := X"00000000";
		ram_buffer(10022) := X"00000000";
		ram_buffer(10023) := X"00000000";
		ram_buffer(10024) := X"00000000";
		ram_buffer(10025) := X"00000000";
		ram_buffer(10026) := X"00000000";
		ram_buffer(10027) := X"00000000";
		ram_buffer(10028) := X"00000000";
		ram_buffer(10029) := X"00000000";
		ram_buffer(10030) := X"00000000";
		ram_buffer(10031) := X"00000000";
		ram_buffer(10032) := X"00000000";
		ram_buffer(10033) := X"00000000";
		ram_buffer(10034) := X"00000000";
		ram_buffer(10035) := X"00000000";
		ram_buffer(10036) := X"00000000";
		ram_buffer(10037) := X"00000000";
		ram_buffer(10038) := X"00000000";
		ram_buffer(10039) := X"00000000";
		ram_buffer(10040) := X"00000000";
		ram_buffer(10041) := X"00000000";
		ram_buffer(10042) := X"00000000";
		ram_buffer(10043) := X"00000000";
		ram_buffer(10044) := X"00000000";
		ram_buffer(10045) := X"00000000";
		ram_buffer(10046) := X"00000000";
		ram_buffer(10047) := X"00000000";
		ram_buffer(10048) := X"00000000";
		ram_buffer(10049) := X"00000000";
		ram_buffer(10050) := X"00000000";
		ram_buffer(10051) := X"00000000";
		ram_buffer(10052) := X"00000000";
		ram_buffer(10053) := X"00000000";
		ram_buffer(10054) := X"00000000";
		ram_buffer(10055) := X"00000000";
		ram_buffer(10056) := X"00000000";
		ram_buffer(10057) := X"00000000";
		ram_buffer(10058) := X"00000000";
		ram_buffer(10059) := X"00000000";
		ram_buffer(10060) := X"00000000";
		ram_buffer(10061) := X"00000000";
		ram_buffer(10062) := X"00000000";
		ram_buffer(10063) := X"00000000";
		ram_buffer(10064) := X"00000000";
		ram_buffer(10065) := X"00000000";
		ram_buffer(10066) := X"00000000";
		ram_buffer(10067) := X"00000000";
		ram_buffer(10068) := X"00000000";
		ram_buffer(10069) := X"00000000";
		ram_buffer(10070) := X"00000000";
		ram_buffer(10071) := X"00000000";
		ram_buffer(10072) := X"00000000";
		ram_buffer(10073) := X"00000000";
		ram_buffer(10074) := X"00000000";
		ram_buffer(10075) := X"00000000";
		ram_buffer(10076) := X"00000000";
		ram_buffer(10077) := X"00000000";
		ram_buffer(10078) := X"00000000";
		ram_buffer(10079) := X"00000000";
		ram_buffer(10080) := X"00000000";
		ram_buffer(10081) := X"00000000";
		ram_buffer(10082) := X"00000000";
		ram_buffer(10083) := X"00000000";
		ram_buffer(10084) := X"00000000";
		ram_buffer(10085) := X"00000000";
		ram_buffer(10086) := X"00000000";
		ram_buffer(10087) := X"00000000";
		ram_buffer(10088) := X"00000000";
		ram_buffer(10089) := X"00000000";
		ram_buffer(10090) := X"00000000";
		ram_buffer(10091) := X"00000000";
		ram_buffer(10092) := X"00000000";
		ram_buffer(10093) := X"00000000";
		ram_buffer(10094) := X"00000000";
		ram_buffer(10095) := X"00000000";
		ram_buffer(10096) := X"00000000";
		ram_buffer(10097) := X"00000000";
		ram_buffer(10098) := X"00000000";
		ram_buffer(10099) := X"00000000";
		ram_buffer(10100) := X"00000000";
		ram_buffer(10101) := X"00000000";
		ram_buffer(10102) := X"00000000";
		ram_buffer(10103) := X"00000000";
		ram_buffer(10104) := X"00000000";
		ram_buffer(10105) := X"00000000";
		ram_buffer(10106) := X"00000000";
		ram_buffer(10107) := X"00000000";
		ram_buffer(10108) := X"00000000";
		ram_buffer(10109) := X"00000000";
		ram_buffer(10110) := X"00000000";
		ram_buffer(10111) := X"00000000";
		ram_buffer(10112) := X"00000000";
		ram_buffer(10113) := X"00000000";
		ram_buffer(10114) := X"00000000";
		ram_buffer(10115) := X"00000000";
		ram_buffer(10116) := X"00000000";
		ram_buffer(10117) := X"00000000";
		ram_buffer(10118) := X"00000000";
		ram_buffer(10119) := X"00000000";
		ram_buffer(10120) := X"00000000";
		ram_buffer(10121) := X"00000000";
		ram_buffer(10122) := X"00000000";
		ram_buffer(10123) := X"00000000";
		ram_buffer(10124) := X"00000000";
		ram_buffer(10125) := X"00000000";
		ram_buffer(10126) := X"00000000";
		ram_buffer(10127) := X"00000000";
		ram_buffer(10128) := X"00000000";
		ram_buffer(10129) := X"00000000";
		ram_buffer(10130) := X"00000000";
		ram_buffer(10131) := X"00000000";
		ram_buffer(10132) := X"00000000";
		ram_buffer(10133) := X"00000000";
		ram_buffer(10134) := X"00000000";
		ram_buffer(10135) := X"00000000";
		ram_buffer(10136) := X"00000000";
		ram_buffer(10137) := X"00000000";
		ram_buffer(10138) := X"00000000";
		ram_buffer(10139) := X"00000000";
		ram_buffer(10140) := X"00000000";
		ram_buffer(10141) := X"00000000";
		ram_buffer(10142) := X"00000000";
		ram_buffer(10143) := X"00000000";
		ram_buffer(10144) := X"00000000";
		ram_buffer(10145) := X"00000000";
		ram_buffer(10146) := X"00000000";
		ram_buffer(10147) := X"00000000";
		ram_buffer(10148) := X"00000000";
		ram_buffer(10149) := X"00000000";
		ram_buffer(10150) := X"00000000";
		ram_buffer(10151) := X"00000000";
		ram_buffer(10152) := X"00000000";
		ram_buffer(10153) := X"00000000";
		ram_buffer(10154) := X"00000000";
		ram_buffer(10155) := X"00000000";
		ram_buffer(10156) := X"00000000";
		ram_buffer(10157) := X"00000000";
		ram_buffer(10158) := X"00000000";
		ram_buffer(10159) := X"00000000";
		ram_buffer(10160) := X"00000000";
		ram_buffer(10161) := X"00000000";
		ram_buffer(10162) := X"00000000";
		ram_buffer(10163) := X"00000000";
		ram_buffer(10164) := X"00000000";
		ram_buffer(10165) := X"00000000";
		ram_buffer(10166) := X"00000000";
		ram_buffer(10167) := X"00000000";
		ram_buffer(10168) := X"00000000";
		ram_buffer(10169) := X"00000000";
		ram_buffer(10170) := X"00000000";
		ram_buffer(10171) := X"00000000";
		ram_buffer(10172) := X"00000000";
		ram_buffer(10173) := X"00000000";
		ram_buffer(10174) := X"00000000";
		ram_buffer(10175) := X"00000000";
		ram_buffer(10176) := X"00000000";
		ram_buffer(10177) := X"00000000";
		ram_buffer(10178) := X"00000000";
		ram_buffer(10179) := X"00000000";
		ram_buffer(10180) := X"00000000";
		ram_buffer(10181) := X"00000000";
		ram_buffer(10182) := X"00000000";
		ram_buffer(10183) := X"00000000";
		ram_buffer(10184) := X"00000000";
		ram_buffer(10185) := X"00000000";
		ram_buffer(10186) := X"00000000";
		ram_buffer(10187) := X"00000000";
		ram_buffer(10188) := X"00000000";
		ram_buffer(10189) := X"00000000";
		ram_buffer(10190) := X"00000000";
		ram_buffer(10191) := X"00000000";
		ram_buffer(10192) := X"00000000";
		ram_buffer(10193) := X"00000000";
		ram_buffer(10194) := X"00000000";
		ram_buffer(10195) := X"00000000";
		ram_buffer(10196) := X"00000000";
		ram_buffer(10197) := X"00000000";
		ram_buffer(10198) := X"00000000";
		ram_buffer(10199) := X"00000000";
		ram_buffer(10200) := X"00000000";
		ram_buffer(10201) := X"00000000";
		ram_buffer(10202) := X"00000000";
		ram_buffer(10203) := X"00000000";
		ram_buffer(10204) := X"00000000";
		ram_buffer(10205) := X"00000000";
		ram_buffer(10206) := X"00000000";
		ram_buffer(10207) := X"00000000";
		ram_buffer(10208) := X"00000000";
		ram_buffer(10209) := X"00000000";
		ram_buffer(10210) := X"00000000";
		ram_buffer(10211) := X"00000000";
		ram_buffer(10212) := X"00000000";
		ram_buffer(10213) := X"00000000";
		ram_buffer(10214) := X"00000000";
		ram_buffer(10215) := X"00000000";
		ram_buffer(10216) := X"00000000";
		ram_buffer(10217) := X"00000000";
		ram_buffer(10218) := X"00000000";
		ram_buffer(10219) := X"00000000";
		ram_buffer(10220) := X"00000000";
		ram_buffer(10221) := X"00000000";
		ram_buffer(10222) := X"00000000";
		ram_buffer(10223) := X"00000000";
		ram_buffer(10224) := X"00000000";
		ram_buffer(10225) := X"00000000";
		ram_buffer(10226) := X"00000000";
		ram_buffer(10227) := X"00000000";
		ram_buffer(10228) := X"00000000";
		ram_buffer(10229) := X"00000000";
		ram_buffer(10230) := X"00000000";
		ram_buffer(10231) := X"00000000";
		ram_buffer(10232) := X"00000000";
		ram_buffer(10233) := X"00000000";
		ram_buffer(10234) := X"00000000";
		ram_buffer(10235) := X"00000000";
		ram_buffer(10236) := X"00000000";
		ram_buffer(10237) := X"00000000";
		ram_buffer(10238) := X"00000000";
		ram_buffer(10239) := X"00000000";
		ram_buffer(10240) := X"00000000";
		ram_buffer(10241) := X"00000000";
		ram_buffer(10242) := X"00000000";
		ram_buffer(10243) := X"00000000";
		ram_buffer(10244) := X"00000000";
		ram_buffer(10245) := X"00000000";
		ram_buffer(10246) := X"00000000";
		ram_buffer(10247) := X"00000000";
		ram_buffer(10248) := X"00000000";
		ram_buffer(10249) := X"00000000";
		ram_buffer(10250) := X"00000000";
		ram_buffer(10251) := X"00000000";
		ram_buffer(10252) := X"00000000";
		ram_buffer(10253) := X"00000000";
		ram_buffer(10254) := X"00000000";
		ram_buffer(10255) := X"00000000";
		ram_buffer(10256) := X"00000000";
		ram_buffer(10257) := X"00000000";
		ram_buffer(10258) := X"00000000";
		ram_buffer(10259) := X"00000000";
		ram_buffer(10260) := X"00000000";
		ram_buffer(10261) := X"00000000";
		ram_buffer(10262) := X"00000000";
		ram_buffer(10263) := X"00000000";
		ram_buffer(10264) := X"00000000";
		ram_buffer(10265) := X"00000000";
		ram_buffer(10266) := X"00000000";
		ram_buffer(10267) := X"00000000";
		ram_buffer(10268) := X"00000000";
		ram_buffer(10269) := X"00000000";
		ram_buffer(10270) := X"00000000";
		ram_buffer(10271) := X"00000000";
		ram_buffer(10272) := X"00000000";
		ram_buffer(10273) := X"00000000";
		ram_buffer(10274) := X"00000000";
		ram_buffer(10275) := X"00000000";
		ram_buffer(10276) := X"00000000";
		ram_buffer(10277) := X"00000000";
		ram_buffer(10278) := X"00000000";
		ram_buffer(10279) := X"00000000";
		ram_buffer(10280) := X"00000000";
		ram_buffer(10281) := X"00000000";
		ram_buffer(10282) := X"00000000";
		ram_buffer(10283) := X"00000000";
		ram_buffer(10284) := X"00000000";
		ram_buffer(10285) := X"00000000";
		ram_buffer(10286) := X"00000000";
		ram_buffer(10287) := X"00000000";
		ram_buffer(10288) := X"00000000";
		ram_buffer(10289) := X"00000000";
		ram_buffer(10290) := X"00000000";
		ram_buffer(10291) := X"00000000";
		ram_buffer(10292) := X"00000000";
		ram_buffer(10293) := X"00000000";
		ram_buffer(10294) := X"00000000";
		ram_buffer(10295) := X"00000000";
		ram_buffer(10296) := X"00000000";
		ram_buffer(10297) := X"00000000";
		ram_buffer(10298) := X"00000000";
		ram_buffer(10299) := X"00000000";
		ram_buffer(10300) := X"00000000";
		ram_buffer(10301) := X"00000000";
		ram_buffer(10302) := X"00000000";
		ram_buffer(10303) := X"00000000";
		ram_buffer(10304) := X"00000000";
		ram_buffer(10305) := X"00000000";
		ram_buffer(10306) := X"00000000";
		ram_buffer(10307) := X"00000000";
		ram_buffer(10308) := X"00000000";
		ram_buffer(10309) := X"00000000";
		ram_buffer(10310) := X"00000000";
		ram_buffer(10311) := X"00000000";
		ram_buffer(10312) := X"00000000";
		ram_buffer(10313) := X"00000000";
		ram_buffer(10314) := X"00000000";
		ram_buffer(10315) := X"00000000";
		ram_buffer(10316) := X"00000000";
		ram_buffer(10317) := X"00000000";
		ram_buffer(10318) := X"00000000";
		ram_buffer(10319) := X"00000000";
		ram_buffer(10320) := X"00000000";
		ram_buffer(10321) := X"00000000";
		ram_buffer(10322) := X"00000000";
		ram_buffer(10323) := X"00000000";
		ram_buffer(10324) := X"00000000";
		ram_buffer(10325) := X"00000000";
		ram_buffer(10326) := X"00000000";
		ram_buffer(10327) := X"00000000";
		ram_buffer(10328) := X"00000000";
		ram_buffer(10329) := X"00000000";
		ram_buffer(10330) := X"00000000";
		ram_buffer(10331) := X"00000000";
		ram_buffer(10332) := X"00000000";
		ram_buffer(10333) := X"00000000";
		ram_buffer(10334) := X"00000000";
		ram_buffer(10335) := X"00000000";
		ram_buffer(10336) := X"00000000";
		ram_buffer(10337) := X"00000000";
		ram_buffer(10338) := X"00000000";
		ram_buffer(10339) := X"00000000";
		ram_buffer(10340) := X"00000000";
		ram_buffer(10341) := X"00000000";
		ram_buffer(10342) := X"00000000";
		ram_buffer(10343) := X"00000000";
		ram_buffer(10344) := X"00000000";
		ram_buffer(10345) := X"00000000";
		ram_buffer(10346) := X"00000000";
		ram_buffer(10347) := X"00000000";
		ram_buffer(10348) := X"00000000";
		ram_buffer(10349) := X"00000000";
		ram_buffer(10350) := X"00000000";
		ram_buffer(10351) := X"00000000";
		ram_buffer(10352) := X"00000000";
		ram_buffer(10353) := X"00000000";
		ram_buffer(10354) := X"00000000";
		ram_buffer(10355) := X"00000000";
		ram_buffer(10356) := X"00000000";
		ram_buffer(10357) := X"00000000";
		ram_buffer(10358) := X"00000000";
		ram_buffer(10359) := X"00000000";
		ram_buffer(10360) := X"00000000";
		ram_buffer(10361) := X"00000000";
		ram_buffer(10362) := X"00000000";
		ram_buffer(10363) := X"00000000";
		ram_buffer(10364) := X"00000000";
		ram_buffer(10365) := X"00000000";
		ram_buffer(10366) := X"00000000";
		ram_buffer(10367) := X"00000000";
		ram_buffer(10368) := X"00000000";
		ram_buffer(10369) := X"00000000";
		ram_buffer(10370) := X"00000000";
		ram_buffer(10371) := X"00000000";
		ram_buffer(10372) := X"00000000";
		ram_buffer(10373) := X"00000000";
		ram_buffer(10374) := X"00000000";
		ram_buffer(10375) := X"00000000";
		ram_buffer(10376) := X"00000000";
		ram_buffer(10377) := X"00000000";
		ram_buffer(10378) := X"00000000";
		ram_buffer(10379) := X"00000000";
		ram_buffer(10380) := X"00000000";
		ram_buffer(10381) := X"00000000";
		ram_buffer(10382) := X"00000000";
		ram_buffer(10383) := X"00000000";
		ram_buffer(10384) := X"00000000";
		ram_buffer(10385) := X"00000000";
		ram_buffer(10386) := X"00000000";
		ram_buffer(10387) := X"00000000";
		ram_buffer(10388) := X"00000000";
		ram_buffer(10389) := X"00000000";
		ram_buffer(10390) := X"00000000";
		ram_buffer(10391) := X"00000000";
		ram_buffer(10392) := X"00000000";
		ram_buffer(10393) := X"00000000";
		ram_buffer(10394) := X"00000000";
		ram_buffer(10395) := X"00000000";
		ram_buffer(10396) := X"00000000";
		ram_buffer(10397) := X"00000000";
		ram_buffer(10398) := X"00000000";
		ram_buffer(10399) := X"00000000";
		ram_buffer(10400) := X"00000000";
		ram_buffer(10401) := X"00000000";
		ram_buffer(10402) := X"00000000";
		ram_buffer(10403) := X"00000000";
		ram_buffer(10404) := X"00000000";
		ram_buffer(10405) := X"00000000";
		ram_buffer(10406) := X"00000000";
		ram_buffer(10407) := X"00000000";
		ram_buffer(10408) := X"00000000";
		ram_buffer(10409) := X"00000000";
		ram_buffer(10410) := X"00000000";
		ram_buffer(10411) := X"00000000";
		ram_buffer(10412) := X"00000000";
		ram_buffer(10413) := X"00000000";
		ram_buffer(10414) := X"00000000";
		ram_buffer(10415) := X"00000000";
		ram_buffer(10416) := X"00000000";
		ram_buffer(10417) := X"00000000";
		ram_buffer(10418) := X"00000000";
		ram_buffer(10419) := X"00000000";
		ram_buffer(10420) := X"00000000";
		ram_buffer(10421) := X"00000000";
		ram_buffer(10422) := X"00000000";
		ram_buffer(10423) := X"00000000";
		ram_buffer(10424) := X"00000000";
		ram_buffer(10425) := X"00000000";
		ram_buffer(10426) := X"00000000";
		ram_buffer(10427) := X"00000000";
		ram_buffer(10428) := X"00000000";
		ram_buffer(10429) := X"00000000";
		ram_buffer(10430) := X"00000000";
		ram_buffer(10431) := X"00000000";
		ram_buffer(10432) := X"00000000";
		ram_buffer(10433) := X"00000000";
		ram_buffer(10434) := X"00000000";
		ram_buffer(10435) := X"00000000";
		ram_buffer(10436) := X"00000000";
		ram_buffer(10437) := X"00000000";
		ram_buffer(10438) := X"00000000";
		ram_buffer(10439) := X"00000000";
		ram_buffer(10440) := X"00000000";
		ram_buffer(10441) := X"00000000";
		ram_buffer(10442) := X"00000000";
		ram_buffer(10443) := X"00000000";
		ram_buffer(10444) := X"00000000";
		ram_buffer(10445) := X"00000000";
		ram_buffer(10446) := X"00000000";
		ram_buffer(10447) := X"00000000";
		ram_buffer(10448) := X"00000000";
		ram_buffer(10449) := X"00000000";
		ram_buffer(10450) := X"00000000";
		ram_buffer(10451) := X"00000000";
		ram_buffer(10452) := X"00000000";
		ram_buffer(10453) := X"00000000";
		ram_buffer(10454) := X"00000000";
		ram_buffer(10455) := X"00000000";
		ram_buffer(10456) := X"00000000";
		ram_buffer(10457) := X"00000000";
		ram_buffer(10458) := X"00000000";
		ram_buffer(10459) := X"00000000";
		ram_buffer(10460) := X"00000000";
		ram_buffer(10461) := X"00000000";
		ram_buffer(10462) := X"00000000";
		ram_buffer(10463) := X"00000000";
		ram_buffer(10464) := X"00000000";
		ram_buffer(10465) := X"00000000";
		ram_buffer(10466) := X"00000000";
		ram_buffer(10467) := X"00000000";
		ram_buffer(10468) := X"00000000";
		ram_buffer(10469) := X"00000000";
		ram_buffer(10470) := X"00000000";
		ram_buffer(10471) := X"00000000";
		ram_buffer(10472) := X"00000000";
		ram_buffer(10473) := X"00000000";
		ram_buffer(10474) := X"00000000";
		ram_buffer(10475) := X"00000000";
		ram_buffer(10476) := X"00000000";
		ram_buffer(10477) := X"00000000";
		ram_buffer(10478) := X"00000000";
		ram_buffer(10479) := X"00000000";
		ram_buffer(10480) := X"00000000";
		ram_buffer(10481) := X"00000000";
		ram_buffer(10482) := X"00000000";
		ram_buffer(10483) := X"00000000";
		ram_buffer(10484) := X"00000000";
		ram_buffer(10485) := X"00000000";
		ram_buffer(10486) := X"00000000";
		ram_buffer(10487) := X"00000000";
		ram_buffer(10488) := X"00000000";
		ram_buffer(10489) := X"00000000";
		ram_buffer(10490) := X"00000000";
		ram_buffer(10491) := X"00000000";
		ram_buffer(10492) := X"00000000";
		ram_buffer(10493) := X"00000000";
		ram_buffer(10494) := X"00000000";
		ram_buffer(10495) := X"00000000";
		ram_buffer(10496) := X"00000000";
		ram_buffer(10497) := X"00000000";
		ram_buffer(10498) := X"00000000";
		ram_buffer(10499) := X"00000000";
		ram_buffer(10500) := X"00000000";
		ram_buffer(10501) := X"00000000";
		ram_buffer(10502) := X"00000000";
		ram_buffer(10503) := X"00000000";
		ram_buffer(10504) := X"00000000";
		ram_buffer(10505) := X"00000000";
		ram_buffer(10506) := X"00000000";
		ram_buffer(10507) := X"00000000";
		ram_buffer(10508) := X"00000000";
		ram_buffer(10509) := X"00000000";
		ram_buffer(10510) := X"00000000";
		ram_buffer(10511) := X"00000000";
		ram_buffer(10512) := X"00000000";
		ram_buffer(10513) := X"00000000";
		ram_buffer(10514) := X"00000000";
		ram_buffer(10515) := X"00000000";
		ram_buffer(10516) := X"00000000";
		ram_buffer(10517) := X"00000000";
		ram_buffer(10518) := X"00000000";
		ram_buffer(10519) := X"00000000";
		ram_buffer(10520) := X"00000000";
		ram_buffer(10521) := X"00000000";
		ram_buffer(10522) := X"00000000";
		ram_buffer(10523) := X"00000000";
		ram_buffer(10524) := X"00000000";
		ram_buffer(10525) := X"00000000";
		ram_buffer(10526) := X"00000000";
		ram_buffer(10527) := X"00000000";
		ram_buffer(10528) := X"00000000";
		ram_buffer(10529) := X"00000000";
		ram_buffer(10530) := X"00000000";
		ram_buffer(10531) := X"00000000";
		ram_buffer(10532) := X"00000000";
		ram_buffer(10533) := X"00000000";
		ram_buffer(10534) := X"00000000";
		ram_buffer(10535) := X"00000000";
		ram_buffer(10536) := X"00000000";
		ram_buffer(10537) := X"00000000";
		ram_buffer(10538) := X"00000000";
		ram_buffer(10539) := X"00000000";
		ram_buffer(10540) := X"00000000";
		ram_buffer(10541) := X"00000000";
		ram_buffer(10542) := X"00000000";
		ram_buffer(10543) := X"00000000";
		ram_buffer(10544) := X"00000000";
		ram_buffer(10545) := X"00000000";
		ram_buffer(10546) := X"00000000";
		ram_buffer(10547) := X"00000000";
		ram_buffer(10548) := X"00000000";
		ram_buffer(10549) := X"00000000";
		ram_buffer(10550) := X"00000000";
		ram_buffer(10551) := X"00000000";
		ram_buffer(10552) := X"00000000";
		ram_buffer(10553) := X"00000000";
		ram_buffer(10554) := X"00000000";
		ram_buffer(10555) := X"00000000";
		ram_buffer(10556) := X"00000000";
		ram_buffer(10557) := X"00000000";
		ram_buffer(10558) := X"00000000";
		ram_buffer(10559) := X"00000000";
		ram_buffer(10560) := X"00000000";
		ram_buffer(10561) := X"00000000";
		ram_buffer(10562) := X"00000000";
		ram_buffer(10563) := X"00000000";
		ram_buffer(10564) := X"00000000";
		ram_buffer(10565) := X"00000000";
		ram_buffer(10566) := X"00000000";
		ram_buffer(10567) := X"00000000";
		ram_buffer(10568) := X"00000000";
		ram_buffer(10569) := X"00000000";
		ram_buffer(10570) := X"00000000";
		ram_buffer(10571) := X"00000000";
		ram_buffer(10572) := X"00000000";
		ram_buffer(10573) := X"00000000";
		ram_buffer(10574) := X"00000000";
		ram_buffer(10575) := X"00000000";
		ram_buffer(10576) := X"00000000";
		ram_buffer(10577) := X"00000000";
		ram_buffer(10578) := X"00000000";
		ram_buffer(10579) := X"00000000";
		ram_buffer(10580) := X"00000000";
		ram_buffer(10581) := X"00000000";
		ram_buffer(10582) := X"00000000";
		ram_buffer(10583) := X"00000000";
		ram_buffer(10584) := X"00000000";
		ram_buffer(10585) := X"00000000";
		ram_buffer(10586) := X"00000000";
		ram_buffer(10587) := X"00000000";
		ram_buffer(10588) := X"00000000";
		ram_buffer(10589) := X"00000000";
		ram_buffer(10590) := X"00000000";
		ram_buffer(10591) := X"00000000";
		ram_buffer(10592) := X"00000000";
		ram_buffer(10593) := X"00000000";
		ram_buffer(10594) := X"00000000";
		ram_buffer(10595) := X"00000000";
		ram_buffer(10596) := X"00000000";
		ram_buffer(10597) := X"00000000";
		ram_buffer(10598) := X"00000000";
		ram_buffer(10599) := X"00000000";
		ram_buffer(10600) := X"00000000";
		ram_buffer(10601) := X"00000000";
		ram_buffer(10602) := X"00000000";
		ram_buffer(10603) := X"00000000";
		ram_buffer(10604) := X"00000000";
		ram_buffer(10605) := X"00000000";
		ram_buffer(10606) := X"00000000";
		ram_buffer(10607) := X"00000000";
		ram_buffer(10608) := X"00000000";
		ram_buffer(10609) := X"00000000";
		ram_buffer(10610) := X"00000000";
		ram_buffer(10611) := X"00000000";
		ram_buffer(10612) := X"00000000";
		ram_buffer(10613) := X"00000000";
		ram_buffer(10614) := X"00000000";
		ram_buffer(10615) := X"00000000";
		ram_buffer(10616) := X"00000000";
		ram_buffer(10617) := X"00000000";
		ram_buffer(10618) := X"00000000";
		ram_buffer(10619) := X"00000000";
		ram_buffer(10620) := X"00000000";
		ram_buffer(10621) := X"00000000";
		ram_buffer(10622) := X"00000000";
		ram_buffer(10623) := X"00000000";
		ram_buffer(10624) := X"00000000";
		ram_buffer(10625) := X"00000000";
		ram_buffer(10626) := X"00000000";
		ram_buffer(10627) := X"00000000";
		ram_buffer(10628) := X"00000000";
		ram_buffer(10629) := X"00000000";
		ram_buffer(10630) := X"00000000";
		ram_buffer(10631) := X"00000000";
		ram_buffer(10632) := X"00000000";
		ram_buffer(10633) := X"00000000";
		ram_buffer(10634) := X"00000000";
		ram_buffer(10635) := X"00000000";
		ram_buffer(10636) := X"00000000";
		ram_buffer(10637) := X"00000000";
		ram_buffer(10638) := X"00000000";
		ram_buffer(10639) := X"00000000";
		ram_buffer(10640) := X"00000000";
		ram_buffer(10641) := X"00000000";
		ram_buffer(10642) := X"00000000";
		ram_buffer(10643) := X"00000000";
		ram_buffer(10644) := X"00000000";
		ram_buffer(10645) := X"00000000";
		ram_buffer(10646) := X"00000000";
		ram_buffer(10647) := X"00000000";
		ram_buffer(10648) := X"00000000";
		ram_buffer(10649) := X"00000000";
		ram_buffer(10650) := X"00000000";
		ram_buffer(10651) := X"00000000";
		ram_buffer(10652) := X"00000000";
		ram_buffer(10653) := X"00000000";
		ram_buffer(10654) := X"00000000";
		ram_buffer(10655) := X"00000000";
		ram_buffer(10656) := X"00000000";
		ram_buffer(10657) := X"00000000";
		ram_buffer(10658) := X"00000000";
		ram_buffer(10659) := X"00000000";
		ram_buffer(10660) := X"00000000";
		ram_buffer(10661) := X"00000000";
		ram_buffer(10662) := X"00000000";
		ram_buffer(10663) := X"00000000";
		ram_buffer(10664) := X"00000000";
		ram_buffer(10665) := X"00000000";
		ram_buffer(10666) := X"00000000";
		ram_buffer(10667) := X"00000000";
		ram_buffer(10668) := X"00000000";
		ram_buffer(10669) := X"00000000";
		ram_buffer(10670) := X"00000000";
		ram_buffer(10671) := X"00000000";
		ram_buffer(10672) := X"00000000";
		ram_buffer(10673) := X"00000000";
		ram_buffer(10674) := X"00000000";
		ram_buffer(10675) := X"00000000";
		ram_buffer(10676) := X"00000000";
		ram_buffer(10677) := X"00000000";
		ram_buffer(10678) := X"00000000";
		ram_buffer(10679) := X"00000000";
		ram_buffer(10680) := X"00000000";
		ram_buffer(10681) := X"00000000";
		ram_buffer(10682) := X"00000000";
		ram_buffer(10683) := X"00000000";
		ram_buffer(10684) := X"00000000";
		ram_buffer(10685) := X"00000000";
		ram_buffer(10686) := X"00000000";
		ram_buffer(10687) := X"00000000";
		ram_buffer(10688) := X"00000000";
		ram_buffer(10689) := X"00000000";
		ram_buffer(10690) := X"00000000";
		ram_buffer(10691) := X"00000000";
		ram_buffer(10692) := X"00000000";
		ram_buffer(10693) := X"00000000";
		ram_buffer(10694) := X"00000000";
		ram_buffer(10695) := X"00000000";
		ram_buffer(10696) := X"00000000";
		ram_buffer(10697) := X"00000000";
		ram_buffer(10698) := X"00000000";
		ram_buffer(10699) := X"00000000";
		ram_buffer(10700) := X"00000000";
		ram_buffer(10701) := X"00000000";
		ram_buffer(10702) := X"00000000";
		ram_buffer(10703) := X"00000000";
		ram_buffer(10704) := X"00000000";
		ram_buffer(10705) := X"00000000";
		ram_buffer(10706) := X"00000000";
		ram_buffer(10707) := X"00000000";
		ram_buffer(10708) := X"00000000";
		ram_buffer(10709) := X"00000000";
		ram_buffer(10710) := X"00000000";
		ram_buffer(10711) := X"00000000";
		ram_buffer(10712) := X"00000000";
		ram_buffer(10713) := X"00000000";
		ram_buffer(10714) := X"00000000";
		ram_buffer(10715) := X"00000000";
		ram_buffer(10716) := X"00000000";
		ram_buffer(10717) := X"00000000";
		ram_buffer(10718) := X"00000000";
		ram_buffer(10719) := X"00000000";
		ram_buffer(10720) := X"00000000";
		ram_buffer(10721) := X"00000000";
		ram_buffer(10722) := X"00000000";
		ram_buffer(10723) := X"00000000";
		ram_buffer(10724) := X"00000000";
		ram_buffer(10725) := X"00000000";
		ram_buffer(10726) := X"00000000";
		ram_buffer(10727) := X"00000000";
		ram_buffer(10728) := X"00000000";
		ram_buffer(10729) := X"00000000";
		ram_buffer(10730) := X"00000000";
		ram_buffer(10731) := X"00000000";
		ram_buffer(10732) := X"00000000";
		ram_buffer(10733) := X"00000000";
		ram_buffer(10734) := X"00000000";
		ram_buffer(10735) := X"00000000";
		ram_buffer(10736) := X"00000000";
		ram_buffer(10737) := X"00000000";
		ram_buffer(10738) := X"00000000";
		ram_buffer(10739) := X"00000000";
		ram_buffer(10740) := X"00000000";
		ram_buffer(10741) := X"00000000";
		ram_buffer(10742) := X"00000000";
		ram_buffer(10743) := X"00000000";
		ram_buffer(10744) := X"00000000";
		ram_buffer(10745) := X"00000000";
		ram_buffer(10746) := X"00000000";
		ram_buffer(10747) := X"00000000";
		ram_buffer(10748) := X"00000000";
		ram_buffer(10749) := X"00000000";
		ram_buffer(10750) := X"00000000";
		ram_buffer(10751) := X"00000000";
		ram_buffer(10752) := X"00000000";
		ram_buffer(10753) := X"00000000";
		ram_buffer(10754) := X"00000000";
		ram_buffer(10755) := X"00000000";
		ram_buffer(10756) := X"00000000";
		ram_buffer(10757) := X"00000000";
		ram_buffer(10758) := X"00000000";
		ram_buffer(10759) := X"00000000";
		ram_buffer(10760) := X"00000000";
		ram_buffer(10761) := X"00000000";
		ram_buffer(10762) := X"00000000";
		ram_buffer(10763) := X"00000000";
		ram_buffer(10764) := X"00000000";
		ram_buffer(10765) := X"00000000";
		ram_buffer(10766) := X"00000000";
		ram_buffer(10767) := X"00000000";
		ram_buffer(10768) := X"00000000";
		ram_buffer(10769) := X"00000000";
		ram_buffer(10770) := X"00000000";
		ram_buffer(10771) := X"00000000";
		ram_buffer(10772) := X"00000000";
		ram_buffer(10773) := X"00000000";
		ram_buffer(10774) := X"00000000";
		ram_buffer(10775) := X"00000000";
		ram_buffer(10776) := X"00000000";
		ram_buffer(10777) := X"00000000";
		ram_buffer(10778) := X"00000000";
		ram_buffer(10779) := X"00000000";
		ram_buffer(10780) := X"00000000";
		ram_buffer(10781) := X"00000000";
		ram_buffer(10782) := X"00000000";
		ram_buffer(10783) := X"00000000";
		ram_buffer(10784) := X"00000000";
		ram_buffer(10785) := X"00000000";
		ram_buffer(10786) := X"00000000";
		ram_buffer(10787) := X"00000000";
		ram_buffer(10788) := X"00000000";
		ram_buffer(10789) := X"00000000";
		ram_buffer(10790) := X"00000000";
		ram_buffer(10791) := X"00000000";
		ram_buffer(10792) := X"00000000";
		ram_buffer(10793) := X"00000000";
		ram_buffer(10794) := X"00000000";
		ram_buffer(10795) := X"00000000";
		ram_buffer(10796) := X"00000000";
		ram_buffer(10797) := X"00000000";
		ram_buffer(10798) := X"00000000";
		ram_buffer(10799) := X"00000000";
		ram_buffer(10800) := X"00000000";
		ram_buffer(10801) := X"00000000";
		ram_buffer(10802) := X"00000000";
		ram_buffer(10803) := X"00000000";
		ram_buffer(10804) := X"00000000";
		ram_buffer(10805) := X"00000000";
		ram_buffer(10806) := X"00000000";
		ram_buffer(10807) := X"00000000";
		ram_buffer(10808) := X"00000000";
		ram_buffer(10809) := X"00000000";
		ram_buffer(10810) := X"00000000";
		ram_buffer(10811) := X"00000000";
		ram_buffer(10812) := X"00000000";
		ram_buffer(10813) := X"00000000";
		ram_buffer(10814) := X"00000000";
		ram_buffer(10815) := X"00000000";
		ram_buffer(10816) := X"00000000";
		ram_buffer(10817) := X"00000000";
		ram_buffer(10818) := X"00000000";
		ram_buffer(10819) := X"00000000";
		ram_buffer(10820) := X"00000000";
		ram_buffer(10821) := X"00000000";
		ram_buffer(10822) := X"00000000";
		ram_buffer(10823) := X"00000000";
		ram_buffer(10824) := X"00000000";
		ram_buffer(10825) := X"00000000";
		ram_buffer(10826) := X"00000000";
		ram_buffer(10827) := X"00000000";
		ram_buffer(10828) := X"00000000";
		ram_buffer(10829) := X"00000000";
		ram_buffer(10830) := X"00000000";
		ram_buffer(10831) := X"00000000";
		ram_buffer(10832) := X"00000000";
		ram_buffer(10833) := X"00000000";
		ram_buffer(10834) := X"00000000";
		ram_buffer(10835) := X"00000000";
		ram_buffer(10836) := X"00000000";
		ram_buffer(10837) := X"00000000";
		ram_buffer(10838) := X"00000000";
		ram_buffer(10839) := X"00000000";
		ram_buffer(10840) := X"00000000";
		ram_buffer(10841) := X"00000000";
		ram_buffer(10842) := X"00000000";
		ram_buffer(10843) := X"00000000";
		ram_buffer(10844) := X"00000000";
		ram_buffer(10845) := X"00000000";
		ram_buffer(10846) := X"00000000";
		ram_buffer(10847) := X"00000000";
		ram_buffer(10848) := X"00000000";
		ram_buffer(10849) := X"00000000";
		ram_buffer(10850) := X"00000000";
		ram_buffer(10851) := X"00000000";
		ram_buffer(10852) := X"00000000";
		ram_buffer(10853) := X"00000000";
		ram_buffer(10854) := X"00000000";
		ram_buffer(10855) := X"00000000";
		ram_buffer(10856) := X"00000000";
		ram_buffer(10857) := X"00000000";
		ram_buffer(10858) := X"00000000";
		ram_buffer(10859) := X"00000000";
		ram_buffer(10860) := X"00000000";
		ram_buffer(10861) := X"00000000";
		ram_buffer(10862) := X"00000000";
		ram_buffer(10863) := X"00000000";
		ram_buffer(10864) := X"00000000";
		ram_buffer(10865) := X"00000000";
		ram_buffer(10866) := X"00000000";
		ram_buffer(10867) := X"00000000";
		ram_buffer(10868) := X"00000000";
		ram_buffer(10869) := X"00000000";
		ram_buffer(10870) := X"00000000";
		ram_buffer(10871) := X"00000000";
		ram_buffer(10872) := X"00000000";
		ram_buffer(10873) := X"00000000";
		ram_buffer(10874) := X"00000000";
		ram_buffer(10875) := X"00000000";
		ram_buffer(10876) := X"00000000";
		ram_buffer(10877) := X"00000000";
		ram_buffer(10878) := X"00000000";
		ram_buffer(10879) := X"00000000";
		ram_buffer(10880) := X"00000000";
		ram_buffer(10881) := X"00000000";
		ram_buffer(10882) := X"00000000";
		ram_buffer(10883) := X"00000000";
		ram_buffer(10884) := X"00000000";
		ram_buffer(10885) := X"00000000";
		ram_buffer(10886) := X"00000000";
		ram_buffer(10887) := X"00000000";
		ram_buffer(10888) := X"00000000";
		ram_buffer(10889) := X"00000000";
		ram_buffer(10890) := X"00000000";
		ram_buffer(10891) := X"00000000";
		ram_buffer(10892) := X"00000000";
		ram_buffer(10893) := X"00000000";
		ram_buffer(10894) := X"00000000";
		ram_buffer(10895) := X"00000000";
		ram_buffer(10896) := X"00000000";
		ram_buffer(10897) := X"00000000";
		ram_buffer(10898) := X"00000000";
		ram_buffer(10899) := X"00000000";
		ram_buffer(10900) := X"00000000";
		ram_buffer(10901) := X"00000000";
		ram_buffer(10902) := X"00000000";
		ram_buffer(10903) := X"00000000";
		ram_buffer(10904) := X"00000000";
		ram_buffer(10905) := X"00000000";
		ram_buffer(10906) := X"00000000";
		ram_buffer(10907) := X"00000000";
		ram_buffer(10908) := X"00000000";
		ram_buffer(10909) := X"00000000";
		ram_buffer(10910) := X"00000000";
		ram_buffer(10911) := X"00000000";
		ram_buffer(10912) := X"00000000";
		ram_buffer(10913) := X"00000000";
		ram_buffer(10914) := X"00000000";
		ram_buffer(10915) := X"00000000";
		ram_buffer(10916) := X"00000000";
		ram_buffer(10917) := X"00000000";
		ram_buffer(10918) := X"00000000";
		ram_buffer(10919) := X"00000000";
		ram_buffer(10920) := X"00000000";
		ram_buffer(10921) := X"00000000";
		ram_buffer(10922) := X"00000000";
		ram_buffer(10923) := X"00000000";
		ram_buffer(10924) := X"00000000";
		ram_buffer(10925) := X"00000000";
		ram_buffer(10926) := X"00000000";
		ram_buffer(10927) := X"00000000";
		ram_buffer(10928) := X"00000000";
		ram_buffer(10929) := X"00000000";
		ram_buffer(10930) := X"00000000";
		ram_buffer(10931) := X"00000000";
		ram_buffer(10932) := X"00000000";
		ram_buffer(10933) := X"00000000";
		ram_buffer(10934) := X"00000000";
		ram_buffer(10935) := X"00000000";
		ram_buffer(10936) := X"00000000";
		ram_buffer(10937) := X"00000000";
		ram_buffer(10938) := X"00000000";
		ram_buffer(10939) := X"00000000";
		ram_buffer(10940) := X"00000000";
		ram_buffer(10941) := X"00000000";
		ram_buffer(10942) := X"00000000";
		ram_buffer(10943) := X"00000000";
		ram_buffer(10944) := X"00000000";
		ram_buffer(10945) := X"00000000";
		ram_buffer(10946) := X"00000000";
		ram_buffer(10947) := X"00000000";
		ram_buffer(10948) := X"00000000";
		ram_buffer(10949) := X"00000000";
		ram_buffer(10950) := X"00000000";
		ram_buffer(10951) := X"00000000";
		ram_buffer(10952) := X"00000000";
		ram_buffer(10953) := X"00000000";
		ram_buffer(10954) := X"00000000";
		ram_buffer(10955) := X"00000000";
		ram_buffer(10956) := X"00000000";
		ram_buffer(10957) := X"00000000";
		ram_buffer(10958) := X"00000000";
		ram_buffer(10959) := X"00000000";
		ram_buffer(10960) := X"00000000";
		ram_buffer(10961) := X"00000000";
		ram_buffer(10962) := X"00000000";
		ram_buffer(10963) := X"00000000";
		ram_buffer(10964) := X"00000000";
		ram_buffer(10965) := X"00000000";
		ram_buffer(10966) := X"00000000";
		ram_buffer(10967) := X"00000000";
		ram_buffer(10968) := X"00000000";
		ram_buffer(10969) := X"00000000";
		ram_buffer(10970) := X"00000000";
		ram_buffer(10971) := X"00000000";
		ram_buffer(10972) := X"00000000";
		ram_buffer(10973) := X"00000000";
		ram_buffer(10974) := X"00000000";
		ram_buffer(10975) := X"00000000";
		ram_buffer(10976) := X"00000000";
		ram_buffer(10977) := X"00000000";
		ram_buffer(10978) := X"00000000";
		ram_buffer(10979) := X"00000000";
		ram_buffer(10980) := X"00000000";
		ram_buffer(10981) := X"00000000";
		ram_buffer(10982) := X"00000000";
		ram_buffer(10983) := X"00000000";
		ram_buffer(10984) := X"00000000";
		ram_buffer(10985) := X"00000000";
		ram_buffer(10986) := X"00000000";
		ram_buffer(10987) := X"00000000";
		ram_buffer(10988) := X"00000000";
		ram_buffer(10989) := X"00000000";
		ram_buffer(10990) := X"00000000";
		ram_buffer(10991) := X"00000000";
		ram_buffer(10992) := X"00000000";
		ram_buffer(10993) := X"00000000";
		ram_buffer(10994) := X"00000000";
		ram_buffer(10995) := X"00000000";
		ram_buffer(10996) := X"00000000";
		ram_buffer(10997) := X"00000000";
		ram_buffer(10998) := X"00000000";
		ram_buffer(10999) := X"00000000";
		ram_buffer(11000) := X"00000000";
		ram_buffer(11001) := X"00000000";
		ram_buffer(11002) := X"00000000";
		ram_buffer(11003) := X"00000000";
		ram_buffer(11004) := X"00000000";
		ram_buffer(11005) := X"00000000";
		ram_buffer(11006) := X"00000000";
		ram_buffer(11007) := X"00000000";
		ram_buffer(11008) := X"00000000";
		ram_buffer(11009) := X"00000000";
		ram_buffer(11010) := X"00000000";
		ram_buffer(11011) := X"00000000";
		ram_buffer(11012) := X"00000000";
		ram_buffer(11013) := X"00000000";
		ram_buffer(11014) := X"00000000";
		ram_buffer(11015) := X"00000000";
		ram_buffer(11016) := X"00000000";
		ram_buffer(11017) := X"00000000";
		ram_buffer(11018) := X"00000000";
		ram_buffer(11019) := X"00000000";
		ram_buffer(11020) := X"00000000";
		ram_buffer(11021) := X"00000000";
		ram_buffer(11022) := X"00000000";
		ram_buffer(11023) := X"00000000";
		ram_buffer(11024) := X"00000000";
		ram_buffer(11025) := X"00000000";
		ram_buffer(11026) := X"00000000";
		ram_buffer(11027) := X"00000000";
		ram_buffer(11028) := X"00000000";
		ram_buffer(11029) := X"00000000";
		ram_buffer(11030) := X"00000000";
		ram_buffer(11031) := X"00000000";
		ram_buffer(11032) := X"00000000";
		ram_buffer(11033) := X"00000000";
		ram_buffer(11034) := X"00000000";
		ram_buffer(11035) := X"00000000";
		ram_buffer(11036) := X"00000000";
		ram_buffer(11037) := X"00000000";
		ram_buffer(11038) := X"00000000";
		ram_buffer(11039) := X"00000000";
		ram_buffer(11040) := X"00000000";
		ram_buffer(11041) := X"00000000";
		ram_buffer(11042) := X"00000000";
		ram_buffer(11043) := X"00000000";
		ram_buffer(11044) := X"00000000";
		ram_buffer(11045) := X"00000000";
		ram_buffer(11046) := X"00000000";
		ram_buffer(11047) := X"00000000";
		ram_buffer(11048) := X"00000000";
		ram_buffer(11049) := X"00000000";
		ram_buffer(11050) := X"00000000";
		ram_buffer(11051) := X"00000000";
		ram_buffer(11052) := X"00000000";
		ram_buffer(11053) := X"00000000";
		ram_buffer(11054) := X"00000000";
		ram_buffer(11055) := X"00000000";
		ram_buffer(11056) := X"00000000";
		ram_buffer(11057) := X"00000000";
		ram_buffer(11058) := X"00000000";
		ram_buffer(11059) := X"00000000";
		ram_buffer(11060) := X"00000000";
		ram_buffer(11061) := X"00000000";
		ram_buffer(11062) := X"00000000";
		ram_buffer(11063) := X"00000000";
		ram_buffer(11064) := X"00000000";
		ram_buffer(11065) := X"00000000";
		ram_buffer(11066) := X"00000000";
		ram_buffer(11067) := X"00000000";
		ram_buffer(11068) := X"00000000";
		ram_buffer(11069) := X"00000000";
		ram_buffer(11070) := X"00000000";
		ram_buffer(11071) := X"00000000";
		ram_buffer(11072) := X"00000000";
		ram_buffer(11073) := X"00000000";
		ram_buffer(11074) := X"00000000";
		ram_buffer(11075) := X"00000000";
		ram_buffer(11076) := X"00000000";
		ram_buffer(11077) := X"00000000";
		ram_buffer(11078) := X"00000000";
		ram_buffer(11079) := X"00000000";
		ram_buffer(11080) := X"00000000";
		ram_buffer(11081) := X"00000000";
		ram_buffer(11082) := X"00000000";
		ram_buffer(11083) := X"00000000";
		ram_buffer(11084) := X"00000000";
		ram_buffer(11085) := X"00000000";
		ram_buffer(11086) := X"00000000";
		ram_buffer(11087) := X"00000000";
		ram_buffer(11088) := X"00000000";
		ram_buffer(11089) := X"00000000";
		ram_buffer(11090) := X"00000000";
		ram_buffer(11091) := X"00000000";
		ram_buffer(11092) := X"00000000";
		ram_buffer(11093) := X"00000000";
		ram_buffer(11094) := X"00000000";
		ram_buffer(11095) := X"00000000";
		ram_buffer(11096) := X"00000000";
		ram_buffer(11097) := X"00000000";
		ram_buffer(11098) := X"00000000";
		ram_buffer(11099) := X"00000000";
		ram_buffer(11100) := X"00000000";
		ram_buffer(11101) := X"00000000";
		ram_buffer(11102) := X"00000000";
		ram_buffer(11103) := X"00000000";
		ram_buffer(11104) := X"00000000";
		ram_buffer(11105) := X"00000000";
		ram_buffer(11106) := X"00000000";
		ram_buffer(11107) := X"00000000";
		ram_buffer(11108) := X"00000000";
		ram_buffer(11109) := X"00000000";
		ram_buffer(11110) := X"00000000";
		ram_buffer(11111) := X"00000000";
		ram_buffer(11112) := X"00000000";
		ram_buffer(11113) := X"00000000";
		ram_buffer(11114) := X"00000000";
		ram_buffer(11115) := X"00000000";
		ram_buffer(11116) := X"00000000";
		ram_buffer(11117) := X"00000000";
		ram_buffer(11118) := X"00000000";
		ram_buffer(11119) := X"00000000";
		ram_buffer(11120) := X"00000000";
		ram_buffer(11121) := X"00000000";
		ram_buffer(11122) := X"00000000";
		ram_buffer(11123) := X"00000000";
		ram_buffer(11124) := X"00000000";
		ram_buffer(11125) := X"00000000";
		ram_buffer(11126) := X"00000000";
		ram_buffer(11127) := X"00000000";
		ram_buffer(11128) := X"00000000";
		ram_buffer(11129) := X"00000000";
		ram_buffer(11130) := X"00000000";
		ram_buffer(11131) := X"00000000";
		ram_buffer(11132) := X"00000000";
		ram_buffer(11133) := X"00000000";
		ram_buffer(11134) := X"00000000";
		ram_buffer(11135) := X"00000000";
		ram_buffer(11136) := X"00000000";
		ram_buffer(11137) := X"00000000";
		ram_buffer(11138) := X"00000000";
		ram_buffer(11139) := X"00000000";
		ram_buffer(11140) := X"00000000";
		ram_buffer(11141) := X"00000000";
		ram_buffer(11142) := X"00000000";
		ram_buffer(11143) := X"00000000";
		ram_buffer(11144) := X"00000000";
		ram_buffer(11145) := X"00000000";
		ram_buffer(11146) := X"00000000";
		ram_buffer(11147) := X"00000000";
		ram_buffer(11148) := X"00000000";
		ram_buffer(11149) := X"00000000";
		ram_buffer(11150) := X"00000000";
		ram_buffer(11151) := X"00000000";
		ram_buffer(11152) := X"00000000";
		ram_buffer(11153) := X"00000000";
		ram_buffer(11154) := X"00000000";
		ram_buffer(11155) := X"00000000";
		ram_buffer(11156) := X"00000000";
		ram_buffer(11157) := X"00000000";
		ram_buffer(11158) := X"00000000";
		ram_buffer(11159) := X"00000000";
		ram_buffer(11160) := X"00000000";
		ram_buffer(11161) := X"00000000";
		ram_buffer(11162) := X"00000000";
		ram_buffer(11163) := X"00000000";
		ram_buffer(11164) := X"00000000";
		ram_buffer(11165) := X"00000000";
		ram_buffer(11166) := X"00000000";
		ram_buffer(11167) := X"00000000";
		ram_buffer(11168) := X"00000000";
		ram_buffer(11169) := X"00000000";
		ram_buffer(11170) := X"00000000";
		ram_buffer(11171) := X"00000000";
		ram_buffer(11172) := X"00000000";
		ram_buffer(11173) := X"00000000";
		ram_buffer(11174) := X"00000000";
		ram_buffer(11175) := X"00000000";
		ram_buffer(11176) := X"00000000";
		ram_buffer(11177) := X"00000000";
		ram_buffer(11178) := X"00000000";
		ram_buffer(11179) := X"00000000";
		ram_buffer(11180) := X"00000000";
		ram_buffer(11181) := X"00000000";
		ram_buffer(11182) := X"00000000";
		ram_buffer(11183) := X"00000000";
		ram_buffer(11184) := X"00000000";
		ram_buffer(11185) := X"00000000";
		ram_buffer(11186) := X"00000000";
		ram_buffer(11187) := X"00000000";
		ram_buffer(11188) := X"00000000";
		ram_buffer(11189) := X"00000000";
		ram_buffer(11190) := X"00000000";
		ram_buffer(11191) := X"00000000";
		ram_buffer(11192) := X"00000000";
		ram_buffer(11193) := X"00000000";
		ram_buffer(11194) := X"00000000";
		ram_buffer(11195) := X"00000000";
		ram_buffer(11196) := X"00000000";
		ram_buffer(11197) := X"00000000";
		ram_buffer(11198) := X"00000000";
		ram_buffer(11199) := X"00000000";
		ram_buffer(11200) := X"00000000";
		ram_buffer(11201) := X"00000000";
		ram_buffer(11202) := X"00000000";
		ram_buffer(11203) := X"00000000";
		ram_buffer(11204) := X"00000000";
		ram_buffer(11205) := X"00000000";
		ram_buffer(11206) := X"00000000";
		ram_buffer(11207) := X"00000000";
		ram_buffer(11208) := X"00000000";
		ram_buffer(11209) := X"00000000";
		ram_buffer(11210) := X"00000000";
		ram_buffer(11211) := X"00000000";
		ram_buffer(11212) := X"00000000";
		ram_buffer(11213) := X"00000000";
		ram_buffer(11214) := X"00000000";
		ram_buffer(11215) := X"00000000";
		ram_buffer(11216) := X"00000000";
		ram_buffer(11217) := X"00000000";
		ram_buffer(11218) := X"00000000";
		ram_buffer(11219) := X"00000000";
		ram_buffer(11220) := X"00000000";
		ram_buffer(11221) := X"00000000";
		ram_buffer(11222) := X"00000000";
		ram_buffer(11223) := X"00000000";
		ram_buffer(11224) := X"00000000";
		ram_buffer(11225) := X"00000000";
		ram_buffer(11226) := X"00000000";
		ram_buffer(11227) := X"00000000";
		ram_buffer(11228) := X"00000000";
		ram_buffer(11229) := X"00000000";
		ram_buffer(11230) := X"00000000";
		ram_buffer(11231) := X"00000000";
		ram_buffer(11232) := X"00000000";
		ram_buffer(11233) := X"00000000";
		ram_buffer(11234) := X"00000000";
		ram_buffer(11235) := X"00000000";
		ram_buffer(11236) := X"00000000";
		ram_buffer(11237) := X"00000000";
		ram_buffer(11238) := X"00000000";
		ram_buffer(11239) := X"00000000";
		ram_buffer(11240) := X"00000000";
		ram_buffer(11241) := X"00000000";
		ram_buffer(11242) := X"00000000";
		ram_buffer(11243) := X"00000000";
		ram_buffer(11244) := X"00000000";
		ram_buffer(11245) := X"00000000";
		ram_buffer(11246) := X"00000000";
		ram_buffer(11247) := X"00000000";
		ram_buffer(11248) := X"00000000";
		ram_buffer(11249) := X"00000000";
		ram_buffer(11250) := X"00000000";
		ram_buffer(11251) := X"00000000";
		ram_buffer(11252) := X"00000000";
		ram_buffer(11253) := X"00000000";
		ram_buffer(11254) := X"00000000";
		ram_buffer(11255) := X"00000000";
		ram_buffer(11256) := X"00000000";
		ram_buffer(11257) := X"00000000";
		ram_buffer(11258) := X"00000000";
		ram_buffer(11259) := X"00000000";
		ram_buffer(11260) := X"00000000";
		ram_buffer(11261) := X"00000000";
		ram_buffer(11262) := X"00000000";
		ram_buffer(11263) := X"00000000";
		ram_buffer(11264) := X"00000000";
		ram_buffer(11265) := X"00000000";
		ram_buffer(11266) := X"00000000";
		ram_buffer(11267) := X"00000000";
		ram_buffer(11268) := X"00000000";
		ram_buffer(11269) := X"00000000";
		ram_buffer(11270) := X"00000000";
		ram_buffer(11271) := X"00000000";
		ram_buffer(11272) := X"00000000";
		ram_buffer(11273) := X"00000000";
		ram_buffer(11274) := X"00000000";
		ram_buffer(11275) := X"00000000";
		ram_buffer(11276) := X"00000000";
		ram_buffer(11277) := X"00000000";
		ram_buffer(11278) := X"00000000";
		ram_buffer(11279) := X"00000000";
		ram_buffer(11280) := X"00000000";
		ram_buffer(11281) := X"00000000";
		ram_buffer(11282) := X"00000000";
		ram_buffer(11283) := X"00000000";
		ram_buffer(11284) := X"00000000";
		ram_buffer(11285) := X"00000000";
		ram_buffer(11286) := X"00000000";
		ram_buffer(11287) := X"00000000";
		ram_buffer(11288) := X"00000000";
		ram_buffer(11289) := X"00000000";
		ram_buffer(11290) := X"00000000";
		ram_buffer(11291) := X"00000000";
		ram_buffer(11292) := X"00000000";
		ram_buffer(11293) := X"00000000";
		ram_buffer(11294) := X"00000000";
		ram_buffer(11295) := X"00000000";
		ram_buffer(11296) := X"00000000";
		ram_buffer(11297) := X"00000000";
		ram_buffer(11298) := X"00000000";
		ram_buffer(11299) := X"00000000";
		ram_buffer(11300) := X"00000000";
		ram_buffer(11301) := X"00000000";
		ram_buffer(11302) := X"00000000";
		ram_buffer(11303) := X"00000000";
		ram_buffer(11304) := X"00000000";
		ram_buffer(11305) := X"00000000";
		ram_buffer(11306) := X"00000000";
		ram_buffer(11307) := X"00000000";
		ram_buffer(11308) := X"00000000";
		ram_buffer(11309) := X"00000000";
		ram_buffer(11310) := X"00000000";
		ram_buffer(11311) := X"00000000";
		ram_buffer(11312) := X"00000000";
		ram_buffer(11313) := X"00000000";
		ram_buffer(11314) := X"00000000";
		ram_buffer(11315) := X"00000000";
		ram_buffer(11316) := X"00000000";
		ram_buffer(11317) := X"00000000";
		ram_buffer(11318) := X"00000000";
		ram_buffer(11319) := X"00000000";
		ram_buffer(11320) := X"00000000";
		ram_buffer(11321) := X"00000000";
		ram_buffer(11322) := X"00000000";
		ram_buffer(11323) := X"00000000";
		ram_buffer(11324) := X"00000000";
		ram_buffer(11325) := X"00000000";
		ram_buffer(11326) := X"00000000";
		ram_buffer(11327) := X"00000000";
		ram_buffer(11328) := X"00000000";
		ram_buffer(11329) := X"00000000";
		ram_buffer(11330) := X"00000000";
		ram_buffer(11331) := X"00000000";
		ram_buffer(11332) := X"00000000";
		ram_buffer(11333) := X"00000000";
		ram_buffer(11334) := X"00000000";
		ram_buffer(11335) := X"00000000";
		ram_buffer(11336) := X"00000000";
		ram_buffer(11337) := X"00000000";
		ram_buffer(11338) := X"00000000";
		ram_buffer(11339) := X"00000000";
		ram_buffer(11340) := X"00000000";
		ram_buffer(11341) := X"00000000";
		ram_buffer(11342) := X"00000000";
		ram_buffer(11343) := X"00000000";
		ram_buffer(11344) := X"00000000";
		ram_buffer(11345) := X"00000000";
		ram_buffer(11346) := X"00000000";
		ram_buffer(11347) := X"00000000";
		ram_buffer(11348) := X"00000000";
		ram_buffer(11349) := X"00000000";
		ram_buffer(11350) := X"00000000";
		ram_buffer(11351) := X"00000000";
		ram_buffer(11352) := X"00000000";
		ram_buffer(11353) := X"00000000";
		ram_buffer(11354) := X"00000000";
		ram_buffer(11355) := X"00000000";
		ram_buffer(11356) := X"00000000";
		ram_buffer(11357) := X"00000000";
		ram_buffer(11358) := X"00000000";
		ram_buffer(11359) := X"00000000";
		ram_buffer(11360) := X"00000000";
		ram_buffer(11361) := X"00000000";
		ram_buffer(11362) := X"00000000";
		ram_buffer(11363) := X"00000000";
		ram_buffer(11364) := X"00000000";
		ram_buffer(11365) := X"00000000";
		ram_buffer(11366) := X"00000000";
		ram_buffer(11367) := X"00000000";
		ram_buffer(11368) := X"00000000";
		ram_buffer(11369) := X"00000000";
		ram_buffer(11370) := X"00000000";
		ram_buffer(11371) := X"00000000";
		ram_buffer(11372) := X"00000000";
		ram_buffer(11373) := X"00000000";
		ram_buffer(11374) := X"00000000";
		ram_buffer(11375) := X"00000000";
		ram_buffer(11376) := X"00000000";
		ram_buffer(11377) := X"00000000";
		ram_buffer(11378) := X"00000000";
		ram_buffer(11379) := X"00000000";
		ram_buffer(11380) := X"00000000";
		ram_buffer(11381) := X"00000000";
		ram_buffer(11382) := X"00000000";
		ram_buffer(11383) := X"00000000";
		ram_buffer(11384) := X"00000000";
		ram_buffer(11385) := X"00000000";
		ram_buffer(11386) := X"00000000";
		ram_buffer(11387) := X"00000000";
		ram_buffer(11388) := X"00000000";
		ram_buffer(11389) := X"00000000";
		ram_buffer(11390) := X"00000000";
		ram_buffer(11391) := X"00000000";
		ram_buffer(11392) := X"00000000";
		ram_buffer(11393) := X"00000000";
		ram_buffer(11394) := X"00000000";
		ram_buffer(11395) := X"00000000";
		ram_buffer(11396) := X"00000000";
		ram_buffer(11397) := X"00000000";
		ram_buffer(11398) := X"00000000";
		ram_buffer(11399) := X"00000000";
		ram_buffer(11400) := X"00000000";
		ram_buffer(11401) := X"00000000";
		ram_buffer(11402) := X"00000000";
		ram_buffer(11403) := X"00000000";
		ram_buffer(11404) := X"00000000";
		ram_buffer(11405) := X"00000000";
		ram_buffer(11406) := X"00000000";
		ram_buffer(11407) := X"00000000";
		ram_buffer(11408) := X"00000000";
		ram_buffer(11409) := X"00000000";
		ram_buffer(11410) := X"00000000";
		ram_buffer(11411) := X"00000000";
		ram_buffer(11412) := X"00000000";
		ram_buffer(11413) := X"00000000";
		ram_buffer(11414) := X"00000000";
		ram_buffer(11415) := X"00000000";
		ram_buffer(11416) := X"00000000";
		ram_buffer(11417) := X"00000000";
		ram_buffer(11418) := X"00000000";
		ram_buffer(11419) := X"00000000";
		ram_buffer(11420) := X"00000000";
		ram_buffer(11421) := X"00000000";
		ram_buffer(11422) := X"00000000";
		ram_buffer(11423) := X"00000000";
		ram_buffer(11424) := X"00000000";
		ram_buffer(11425) := X"00000000";
		ram_buffer(11426) := X"00000000";
		ram_buffer(11427) := X"00000000";
		ram_buffer(11428) := X"00000000";
		ram_buffer(11429) := X"00000000";
		ram_buffer(11430) := X"00000000";
		ram_buffer(11431) := X"00000000";
		ram_buffer(11432) := X"00000000";
		ram_buffer(11433) := X"00000000";
		ram_buffer(11434) := X"00000000";
		ram_buffer(11435) := X"00000000";
		ram_buffer(11436) := X"00000000";
		ram_buffer(11437) := X"00000000";
		ram_buffer(11438) := X"00000000";
		ram_buffer(11439) := X"00000000";
		ram_buffer(11440) := X"00000000";
		ram_buffer(11441) := X"00000000";
		ram_buffer(11442) := X"00000000";
		ram_buffer(11443) := X"00000000";
		ram_buffer(11444) := X"00000000";
		ram_buffer(11445) := X"00000000";
		ram_buffer(11446) := X"00000000";
		ram_buffer(11447) := X"00000000";
		ram_buffer(11448) := X"00000000";
		ram_buffer(11449) := X"00000000";
		ram_buffer(11450) := X"00000000";
		ram_buffer(11451) := X"00000000";
		ram_buffer(11452) := X"00000000";
		ram_buffer(11453) := X"00000000";
		ram_buffer(11454) := X"00000000";
		ram_buffer(11455) := X"00000000";
		ram_buffer(11456) := X"00000000";
		ram_buffer(11457) := X"00000000";
		ram_buffer(11458) := X"00000000";
		ram_buffer(11459) := X"00000000";
		ram_buffer(11460) := X"00000000";
		ram_buffer(11461) := X"00000000";
		ram_buffer(11462) := X"00000000";
		ram_buffer(11463) := X"00000000";
		ram_buffer(11464) := X"00000000";
		ram_buffer(11465) := X"00000000";
		ram_buffer(11466) := X"00000000";
		ram_buffer(11467) := X"00000000";
		ram_buffer(11468) := X"00000000";
		ram_buffer(11469) := X"00000000";
		ram_buffer(11470) := X"00000000";
		ram_buffer(11471) := X"00000000";
		ram_buffer(11472) := X"00000000";
		ram_buffer(11473) := X"00000000";
		ram_buffer(11474) := X"00000000";
		ram_buffer(11475) := X"00000000";
		ram_buffer(11476) := X"00000000";
		ram_buffer(11477) := X"00000000";
		ram_buffer(11478) := X"00000000";
		ram_buffer(11479) := X"00000000";
		ram_buffer(11480) := X"00000000";
		ram_buffer(11481) := X"00000000";
		ram_buffer(11482) := X"00000000";
		ram_buffer(11483) := X"00000000";
		ram_buffer(11484) := X"00000000";
		ram_buffer(11485) := X"00000000";
		ram_buffer(11486) := X"00000000";
		ram_buffer(11487) := X"00000000";
		ram_buffer(11488) := X"00000000";
		ram_buffer(11489) := X"00000000";
		ram_buffer(11490) := X"00000000";
		ram_buffer(11491) := X"00000000";
		ram_buffer(11492) := X"00000000";
		ram_buffer(11493) := X"00000000";
		ram_buffer(11494) := X"00000000";
		ram_buffer(11495) := X"00000000";
		ram_buffer(11496) := X"00000000";
		ram_buffer(11497) := X"00000000";
		ram_buffer(11498) := X"00000000";
		ram_buffer(11499) := X"00000000";
		ram_buffer(11500) := X"00000000";
		ram_buffer(11501) := X"00000000";
		ram_buffer(11502) := X"00000000";
		ram_buffer(11503) := X"00000000";
		ram_buffer(11504) := X"00000000";
		ram_buffer(11505) := X"00000000";
		ram_buffer(11506) := X"00000000";
		ram_buffer(11507) := X"00000000";
		ram_buffer(11508) := X"00000000";
		ram_buffer(11509) := X"00000000";
		ram_buffer(11510) := X"00000000";
		ram_buffer(11511) := X"00000000";
		ram_buffer(11512) := X"00000000";
		ram_buffer(11513) := X"00000000";
		ram_buffer(11514) := X"00000000";
		ram_buffer(11515) := X"00000000";
		ram_buffer(11516) := X"00000000";
		ram_buffer(11517) := X"00000000";
		ram_buffer(11518) := X"00000000";
		ram_buffer(11519) := X"00000000";
		ram_buffer(11520) := X"00000000";
		ram_buffer(11521) := X"00000000";
		ram_buffer(11522) := X"00000000";
		ram_buffer(11523) := X"00000000";
		ram_buffer(11524) := X"00000000";
		ram_buffer(11525) := X"00000000";
		ram_buffer(11526) := X"00000000";
		ram_buffer(11527) := X"00000000";
		ram_buffer(11528) := X"00000000";
		ram_buffer(11529) := X"00000000";
		ram_buffer(11530) := X"00000000";
		ram_buffer(11531) := X"00000000";
		ram_buffer(11532) := X"00000000";
		ram_buffer(11533) := X"00000000";
		ram_buffer(11534) := X"00000000";
		ram_buffer(11535) := X"00000000";
		ram_buffer(11536) := X"00000000";
		ram_buffer(11537) := X"00000000";
		ram_buffer(11538) := X"00000000";
		ram_buffer(11539) := X"00000000";
		ram_buffer(11540) := X"00000000";
		ram_buffer(11541) := X"00000000";
		ram_buffer(11542) := X"00000000";
		ram_buffer(11543) := X"00000000";
		ram_buffer(11544) := X"00000000";
		ram_buffer(11545) := X"00000000";
		ram_buffer(11546) := X"00000000";
		ram_buffer(11547) := X"00000000";
		ram_buffer(11548) := X"00000000";
		ram_buffer(11549) := X"00000000";
		ram_buffer(11550) := X"00000000";
		ram_buffer(11551) := X"00000000";
		ram_buffer(11552) := X"00000000";
		ram_buffer(11553) := X"00000000";
		ram_buffer(11554) := X"00000000";
		ram_buffer(11555) := X"00000000";
		ram_buffer(11556) := X"00000000";
		ram_buffer(11557) := X"00000000";
		ram_buffer(11558) := X"00000000";
		ram_buffer(11559) := X"00000000";
		ram_buffer(11560) := X"00000000";
		ram_buffer(11561) := X"00000000";
		ram_buffer(11562) := X"00000000";
		ram_buffer(11563) := X"00000000";
		ram_buffer(11564) := X"00000000";
		ram_buffer(11565) := X"00000000";
		ram_buffer(11566) := X"00000000";
		ram_buffer(11567) := X"00000000";
		ram_buffer(11568) := X"00000000";
		ram_buffer(11569) := X"00000000";
		ram_buffer(11570) := X"00000000";
		ram_buffer(11571) := X"00000000";
		ram_buffer(11572) := X"00000000";
		ram_buffer(11573) := X"00000000";
		ram_buffer(11574) := X"00000000";
		ram_buffer(11575) := X"00000000";
		ram_buffer(11576) := X"00000000";
		ram_buffer(11577) := X"00000000";
		ram_buffer(11578) := X"00000000";
		ram_buffer(11579) := X"00000000";
		ram_buffer(11580) := X"00000000";
		ram_buffer(11581) := X"00000000";
		ram_buffer(11582) := X"00000000";
		ram_buffer(11583) := X"00000000";
		ram_buffer(11584) := X"00000000";
		ram_buffer(11585) := X"00000000";
		ram_buffer(11586) := X"00000000";
		ram_buffer(11587) := X"00000000";
		ram_buffer(11588) := X"00000000";
		ram_buffer(11589) := X"00000000";
		ram_buffer(11590) := X"00000000";
		ram_buffer(11591) := X"00000000";
		ram_buffer(11592) := X"00000000";
		ram_buffer(11593) := X"00000000";
		ram_buffer(11594) := X"00000000";
		ram_buffer(11595) := X"00000000";
		ram_buffer(11596) := X"00000000";
		ram_buffer(11597) := X"00000000";
		ram_buffer(11598) := X"00000000";
		ram_buffer(11599) := X"00000000";
		ram_buffer(11600) := X"00000000";
		ram_buffer(11601) := X"00000000";
		ram_buffer(11602) := X"00000000";
		ram_buffer(11603) := X"00000000";
		ram_buffer(11604) := X"00000000";
		ram_buffer(11605) := X"00000000";
		ram_buffer(11606) := X"00000000";
		ram_buffer(11607) := X"00000000";
		ram_buffer(11608) := X"00000000";
		ram_buffer(11609) := X"00000000";
		ram_buffer(11610) := X"00000000";
		ram_buffer(11611) := X"00000000";
		ram_buffer(11612) := X"00000000";
		ram_buffer(11613) := X"00000000";
		ram_buffer(11614) := X"00000000";
		ram_buffer(11615) := X"00000000";
		ram_buffer(11616) := X"00000000";
		ram_buffer(11617) := X"00000000";
		ram_buffer(11618) := X"00000000";
		ram_buffer(11619) := X"00000000";
		ram_buffer(11620) := X"00000000";
		ram_buffer(11621) := X"00000000";
		ram_buffer(11622) := X"00000000";
		ram_buffer(11623) := X"00000000";
		ram_buffer(11624) := X"00000000";
		ram_buffer(11625) := X"00000000";
		ram_buffer(11626) := X"00000000";
		ram_buffer(11627) := X"00000000";
		ram_buffer(11628) := X"00000000";
		ram_buffer(11629) := X"00000000";
		ram_buffer(11630) := X"00000000";
		ram_buffer(11631) := X"00000000";
		ram_buffer(11632) := X"00000000";
		ram_buffer(11633) := X"00000000";
		ram_buffer(11634) := X"00000000";
		ram_buffer(11635) := X"00000000";
		ram_buffer(11636) := X"00000000";
		ram_buffer(11637) := X"00000000";
		ram_buffer(11638) := X"00000000";
		ram_buffer(11639) := X"00000000";
		ram_buffer(11640) := X"00000000";
		ram_buffer(11641) := X"00000000";
		ram_buffer(11642) := X"00000000";
		ram_buffer(11643) := X"00000000";
		ram_buffer(11644) := X"00000000";
		ram_buffer(11645) := X"00000000";
		ram_buffer(11646) := X"00000000";
		ram_buffer(11647) := X"00000000";
		ram_buffer(11648) := X"00000000";
		ram_buffer(11649) := X"00000000";
		ram_buffer(11650) := X"00000000";
		ram_buffer(11651) := X"00000000";
		ram_buffer(11652) := X"00000000";
		ram_buffer(11653) := X"00000000";
		ram_buffer(11654) := X"00000000";
		ram_buffer(11655) := X"00000000";
		ram_buffer(11656) := X"00000000";
		ram_buffer(11657) := X"00000000";
		ram_buffer(11658) := X"00000000";
		ram_buffer(11659) := X"00000000";
		ram_buffer(11660) := X"00000000";
		ram_buffer(11661) := X"00000000";
		ram_buffer(11662) := X"00000000";
		ram_buffer(11663) := X"00000000";
		ram_buffer(11664) := X"00000000";
		ram_buffer(11665) := X"00000000";
		ram_buffer(11666) := X"00000000";
		ram_buffer(11667) := X"00000000";
		ram_buffer(11668) := X"00000000";
		ram_buffer(11669) := X"00000000";
		ram_buffer(11670) := X"00000000";
		ram_buffer(11671) := X"00000000";
		ram_buffer(11672) := X"00000000";
		ram_buffer(11673) := X"00000000";
		ram_buffer(11674) := X"00000000";
		ram_buffer(11675) := X"00000000";
		ram_buffer(11676) := X"00000000";
		ram_buffer(11677) := X"00000000";
		ram_buffer(11678) := X"00000000";
		ram_buffer(11679) := X"00000000";
		ram_buffer(11680) := X"00000000";
		ram_buffer(11681) := X"00000000";
		ram_buffer(11682) := X"00000000";
		ram_buffer(11683) := X"00000000";
		ram_buffer(11684) := X"00000000";
		ram_buffer(11685) := X"00000000";
		ram_buffer(11686) := X"00000000";
		ram_buffer(11687) := X"00000000";
		ram_buffer(11688) := X"00000000";
		ram_buffer(11689) := X"00000000";
		ram_buffer(11690) := X"00000000";
		ram_buffer(11691) := X"00000000";
		ram_buffer(11692) := X"00000000";
		ram_buffer(11693) := X"00000000";
		ram_buffer(11694) := X"00000000";
		ram_buffer(11695) := X"00000000";
		ram_buffer(11696) := X"00000000";
		ram_buffer(11697) := X"00000000";
		ram_buffer(11698) := X"00000000";
		ram_buffer(11699) := X"00000000";
		ram_buffer(11700) := X"00000000";
		ram_buffer(11701) := X"00000000";
		ram_buffer(11702) := X"00000000";
		ram_buffer(11703) := X"00000000";
		ram_buffer(11704) := X"00000000";
		ram_buffer(11705) := X"00000000";
		ram_buffer(11706) := X"00000000";
		ram_buffer(11707) := X"00000000";
		ram_buffer(11708) := X"00000000";
		ram_buffer(11709) := X"00000000";
		ram_buffer(11710) := X"00000000";
		ram_buffer(11711) := X"00000000";
		ram_buffer(11712) := X"00000000";
		ram_buffer(11713) := X"00000000";
		ram_buffer(11714) := X"00000000";
		ram_buffer(11715) := X"00000000";
		ram_buffer(11716) := X"00000000";
		ram_buffer(11717) := X"00000000";
		ram_buffer(11718) := X"00000000";
		ram_buffer(11719) := X"00000000";
		ram_buffer(11720) := X"00000000";
		ram_buffer(11721) := X"00000000";
		ram_buffer(11722) := X"00000000";
		ram_buffer(11723) := X"00000000";
		ram_buffer(11724) := X"00000000";
		ram_buffer(11725) := X"00000000";
		ram_buffer(11726) := X"00000000";
		ram_buffer(11727) := X"00000000";
		ram_buffer(11728) := X"00000000";
		ram_buffer(11729) := X"00000000";
		ram_buffer(11730) := X"00000000";
		ram_buffer(11731) := X"00000000";
		ram_buffer(11732) := X"00000000";
		ram_buffer(11733) := X"00000000";
		ram_buffer(11734) := X"00000000";
		ram_buffer(11735) := X"00000000";
		ram_buffer(11736) := X"00000000";
		ram_buffer(11737) := X"00000000";
		ram_buffer(11738) := X"00000000";
		ram_buffer(11739) := X"00000000";
		ram_buffer(11740) := X"00000000";
		ram_buffer(11741) := X"00000000";
		ram_buffer(11742) := X"00000000";
		ram_buffer(11743) := X"00000000";
		ram_buffer(11744) := X"00000000";
		ram_buffer(11745) := X"00000000";
		ram_buffer(11746) := X"00000000";
		ram_buffer(11747) := X"00000000";
		ram_buffer(11748) := X"00000000";
		ram_buffer(11749) := X"00000000";
		ram_buffer(11750) := X"00000000";
		ram_buffer(11751) := X"00000000";
		ram_buffer(11752) := X"00000000";
		ram_buffer(11753) := X"00000000";
		ram_buffer(11754) := X"00000000";
		ram_buffer(11755) := X"00000000";
		ram_buffer(11756) := X"00000000";
		ram_buffer(11757) := X"00000000";
		ram_buffer(11758) := X"00000000";
		ram_buffer(11759) := X"00000000";
		ram_buffer(11760) := X"00000000";
		ram_buffer(11761) := X"00000000";
		ram_buffer(11762) := X"00000000";
		ram_buffer(11763) := X"00000000";
		ram_buffer(11764) := X"00000000";
		ram_buffer(11765) := X"00000000";
		ram_buffer(11766) := X"00000000";
		ram_buffer(11767) := X"00000000";
		ram_buffer(11768) := X"00000000";
		ram_buffer(11769) := X"00000000";
		ram_buffer(11770) := X"00000000";
		ram_buffer(11771) := X"00000000";
		ram_buffer(11772) := X"00000000";
		ram_buffer(11773) := X"00000000";
		ram_buffer(11774) := X"00000000";
		ram_buffer(11775) := X"00000000";
		ram_buffer(11776) := X"00000000";
		ram_buffer(11777) := X"00000000";
		ram_buffer(11778) := X"00000000";
		ram_buffer(11779) := X"00000000";
		ram_buffer(11780) := X"00000000";
		ram_buffer(11781) := X"00000000";
		ram_buffer(11782) := X"00000000";
		ram_buffer(11783) := X"00000000";
		ram_buffer(11784) := X"00000000";
		ram_buffer(11785) := X"00000000";
		ram_buffer(11786) := X"00000000";
		ram_buffer(11787) := X"00000000";
		ram_buffer(11788) := X"00000000";
		ram_buffer(11789) := X"00000000";
		ram_buffer(11790) := X"00000000";
		ram_buffer(11791) := X"00000000";
		ram_buffer(11792) := X"00000000";
		ram_buffer(11793) := X"00000000";
		ram_buffer(11794) := X"00000000";
		ram_buffer(11795) := X"00000000";
		ram_buffer(11796) := X"00000000";
		ram_buffer(11797) := X"00000000";
		ram_buffer(11798) := X"00000000";
		ram_buffer(11799) := X"00000000";
		ram_buffer(11800) := X"00000000";
		ram_buffer(11801) := X"00000000";
		ram_buffer(11802) := X"00000000";
		ram_buffer(11803) := X"00000000";
		ram_buffer(11804) := X"00000000";
		ram_buffer(11805) := X"00000000";
		ram_buffer(11806) := X"00000000";
		ram_buffer(11807) := X"00000000";
		ram_buffer(11808) := X"00000000";
		ram_buffer(11809) := X"00000000";
		ram_buffer(11810) := X"00000000";
		ram_buffer(11811) := X"00000000";
		ram_buffer(11812) := X"00000000";
		ram_buffer(11813) := X"00000000";
		ram_buffer(11814) := X"00000000";
		ram_buffer(11815) := X"00000000";
		ram_buffer(11816) := X"00000000";
		ram_buffer(11817) := X"00000000";
		ram_buffer(11818) := X"00000000";
		ram_buffer(11819) := X"00000000";
		ram_buffer(11820) := X"00000000";
		ram_buffer(11821) := X"00000000";
		ram_buffer(11822) := X"00000000";
		ram_buffer(11823) := X"00000000";
		ram_buffer(11824) := X"00000000";
		ram_buffer(11825) := X"00000000";
		ram_buffer(11826) := X"00000000";
		ram_buffer(11827) := X"00000000";
		ram_buffer(11828) := X"00000000";
		ram_buffer(11829) := X"00000000";
		ram_buffer(11830) := X"00000000";
		ram_buffer(11831) := X"00000000";
		ram_buffer(11832) := X"00000000";
		ram_buffer(11833) := X"00000000";
		ram_buffer(11834) := X"00000000";
		ram_buffer(11835) := X"00000000";
		ram_buffer(11836) := X"00000000";
		ram_buffer(11837) := X"00000000";
		ram_buffer(11838) := X"00000000";
		ram_buffer(11839) := X"00000000";
		ram_buffer(11840) := X"00000000";
		ram_buffer(11841) := X"00000000";
		ram_buffer(11842) := X"00000000";
		ram_buffer(11843) := X"00000000";
		ram_buffer(11844) := X"00000000";
		ram_buffer(11845) := X"00000000";
		ram_buffer(11846) := X"00000000";
		ram_buffer(11847) := X"00000000";
		ram_buffer(11848) := X"00000000";
		ram_buffer(11849) := X"00000000";
		ram_buffer(11850) := X"00000000";
		ram_buffer(11851) := X"00000000";
		ram_buffer(11852) := X"00000000";
		ram_buffer(11853) := X"00000000";
		ram_buffer(11854) := X"00000000";
		ram_buffer(11855) := X"00000000";
		ram_buffer(11856) := X"00000000";
		ram_buffer(11857) := X"00000000";
		ram_buffer(11858) := X"00000000";
		ram_buffer(11859) := X"00000000";
		ram_buffer(11860) := X"00000000";
		ram_buffer(11861) := X"00000000";
		ram_buffer(11862) := X"00000000";
		ram_buffer(11863) := X"00000000";
		ram_buffer(11864) := X"00000000";
		ram_buffer(11865) := X"00000000";
		ram_buffer(11866) := X"00000000";
		ram_buffer(11867) := X"00000000";
		ram_buffer(11868) := X"00000000";
		ram_buffer(11869) := X"00000000";
		ram_buffer(11870) := X"00000000";
		ram_buffer(11871) := X"00000000";
		ram_buffer(11872) := X"00000000";
		ram_buffer(11873) := X"00000000";
		ram_buffer(11874) := X"00000000";
		ram_buffer(11875) := X"00000000";
		ram_buffer(11876) := X"00000000";
		ram_buffer(11877) := X"00000000";
		ram_buffer(11878) := X"00000000";
		ram_buffer(11879) := X"00000000";
		ram_buffer(11880) := X"00000000";
		ram_buffer(11881) := X"00000000";
		ram_buffer(11882) := X"00000000";
		ram_buffer(11883) := X"00000000";
		ram_buffer(11884) := X"00000000";
		ram_buffer(11885) := X"00000000";
		ram_buffer(11886) := X"00000000";
		ram_buffer(11887) := X"00000000";
		ram_buffer(11888) := X"00000000";
		ram_buffer(11889) := X"00000000";
		ram_buffer(11890) := X"00000000";
		ram_buffer(11891) := X"00000000";
		ram_buffer(11892) := X"00000000";
		ram_buffer(11893) := X"00000000";
		ram_buffer(11894) := X"00000000";
		ram_buffer(11895) := X"00000000";
		ram_buffer(11896) := X"00000000";
		ram_buffer(11897) := X"00000000";
		ram_buffer(11898) := X"00000000";
		ram_buffer(11899) := X"00000000";
		ram_buffer(11900) := X"00000000";
		ram_buffer(11901) := X"00000000";
		ram_buffer(11902) := X"00000000";
		ram_buffer(11903) := X"00000000";
		ram_buffer(11904) := X"00000000";
		ram_buffer(11905) := X"00000000";
		ram_buffer(11906) := X"00000000";
		ram_buffer(11907) := X"00000000";
		ram_buffer(11908) := X"00000000";
		ram_buffer(11909) := X"00000000";
		ram_buffer(11910) := X"00000000";
		ram_buffer(11911) := X"00000000";
		ram_buffer(11912) := X"00000000";
		ram_buffer(11913) := X"00000000";
		ram_buffer(11914) := X"00000000";
		ram_buffer(11915) := X"00000000";
		ram_buffer(11916) := X"00000000";
		ram_buffer(11917) := X"00000000";
		ram_buffer(11918) := X"00000000";
		ram_buffer(11919) := X"00000000";
		ram_buffer(11920) := X"00000000";
		ram_buffer(11921) := X"00000000";
		ram_buffer(11922) := X"00000000";
		ram_buffer(11923) := X"00000000";
		ram_buffer(11924) := X"00000000";
		ram_buffer(11925) := X"00000000";
		ram_buffer(11926) := X"00000000";
		ram_buffer(11927) := X"00000000";
		ram_buffer(11928) := X"00000000";
		ram_buffer(11929) := X"00000000";
		ram_buffer(11930) := X"00000000";
		ram_buffer(11931) := X"00000000";
		ram_buffer(11932) := X"00000000";
		ram_buffer(11933) := X"00000000";
		ram_buffer(11934) := X"00000000";
		ram_buffer(11935) := X"00000000";
		ram_buffer(11936) := X"00000000";
		ram_buffer(11937) := X"00000000";
		ram_buffer(11938) := X"00000000";
		ram_buffer(11939) := X"00000000";
		ram_buffer(11940) := X"00000000";
		ram_buffer(11941) := X"00000000";
		ram_buffer(11942) := X"00000000";
		ram_buffer(11943) := X"00000000";
		ram_buffer(11944) := X"00000000";
		ram_buffer(11945) := X"00000000";
		ram_buffer(11946) := X"00000000";
		ram_buffer(11947) := X"00000000";
		ram_buffer(11948) := X"00000000";
		ram_buffer(11949) := X"00000000";
		ram_buffer(11950) := X"00000000";
		ram_buffer(11951) := X"00000000";
		ram_buffer(11952) := X"00000000";
		ram_buffer(11953) := X"00000000";
		ram_buffer(11954) := X"00000000";
		ram_buffer(11955) := X"00000000";
		ram_buffer(11956) := X"00000000";
		ram_buffer(11957) := X"00000000";
		ram_buffer(11958) := X"00000000";
		ram_buffer(11959) := X"00000000";
		ram_buffer(11960) := X"00000000";
		ram_buffer(11961) := X"00000000";
		ram_buffer(11962) := X"00000000";
		ram_buffer(11963) := X"00000000";
		ram_buffer(11964) := X"00000000";
		ram_buffer(11965) := X"00000000";
		ram_buffer(11966) := X"00000000";
		ram_buffer(11967) := X"00000000";
		ram_buffer(11968) := X"00000000";
		ram_buffer(11969) := X"00000000";
		ram_buffer(11970) := X"00000000";
		ram_buffer(11971) := X"00000000";
		ram_buffer(11972) := X"00000000";
		ram_buffer(11973) := X"00000000";
		ram_buffer(11974) := X"00000000";
		ram_buffer(11975) := X"00000000";
		ram_buffer(11976) := X"00000000";
		ram_buffer(11977) := X"00000000";
		ram_buffer(11978) := X"00000000";
		ram_buffer(11979) := X"00000000";
		ram_buffer(11980) := X"00000000";
		ram_buffer(11981) := X"00000000";
		ram_buffer(11982) := X"00000000";
		ram_buffer(11983) := X"00000000";
		ram_buffer(11984) := X"00000000";
		ram_buffer(11985) := X"00000000";
		ram_buffer(11986) := X"00000000";
		ram_buffer(11987) := X"00000000";
		ram_buffer(11988) := X"00000000";
		ram_buffer(11989) := X"00000000";
		ram_buffer(11990) := X"00000000";
		ram_buffer(11991) := X"00000000";
		ram_buffer(11992) := X"00000000";
		ram_buffer(11993) := X"00000000";
		ram_buffer(11994) := X"00000000";
		ram_buffer(11995) := X"00000000";
		ram_buffer(11996) := X"00000000";
		ram_buffer(11997) := X"00000000";
		ram_buffer(11998) := X"00000000";
		ram_buffer(11999) := X"00000000";
		ram_buffer(12000) := X"00000000";
		ram_buffer(12001) := X"00000000";
		ram_buffer(12002) := X"00000000";
		ram_buffer(12003) := X"00000000";
		ram_buffer(12004) := X"00000000";
		ram_buffer(12005) := X"00000000";
		ram_buffer(12006) := X"00000000";
		ram_buffer(12007) := X"00000000";
		ram_buffer(12008) := X"00000000";
		ram_buffer(12009) := X"00000000";
		ram_buffer(12010) := X"00000000";
		ram_buffer(12011) := X"00000000";
		ram_buffer(12012) := X"00000000";
		ram_buffer(12013) := X"00000000";
		ram_buffer(12014) := X"00000000";
		ram_buffer(12015) := X"00000000";
		ram_buffer(12016) := X"00000000";
		ram_buffer(12017) := X"00000000";
		ram_buffer(12018) := X"00000000";
		ram_buffer(12019) := X"00000000";
		ram_buffer(12020) := X"00000000";
		ram_buffer(12021) := X"00000000";
		ram_buffer(12022) := X"00000000";
		ram_buffer(12023) := X"00000000";
		ram_buffer(12024) := X"00000000";
		ram_buffer(12025) := X"00000000";
		ram_buffer(12026) := X"00000000";
		ram_buffer(12027) := X"00000000";
		ram_buffer(12028) := X"00000000";
		ram_buffer(12029) := X"00000000";
		ram_buffer(12030) := X"00000000";
		ram_buffer(12031) := X"00000000";
		ram_buffer(12032) := X"00000000";
		ram_buffer(12033) := X"00000000";
		ram_buffer(12034) := X"00000000";
		ram_buffer(12035) := X"00000000";
		ram_buffer(12036) := X"00000000";
		ram_buffer(12037) := X"00000000";
		ram_buffer(12038) := X"00000000";
		ram_buffer(12039) := X"00000000";
		ram_buffer(12040) := X"00000000";
		ram_buffer(12041) := X"00000000";
		ram_buffer(12042) := X"00000000";
		ram_buffer(12043) := X"00000000";
		ram_buffer(12044) := X"00000000";
		ram_buffer(12045) := X"00000000";
		ram_buffer(12046) := X"00000000";
		ram_buffer(12047) := X"00000000";
		ram_buffer(12048) := X"00000000";
		ram_buffer(12049) := X"00000000";
		ram_buffer(12050) := X"00000000";
		ram_buffer(12051) := X"00000000";
		ram_buffer(12052) := X"00000000";
		ram_buffer(12053) := X"00000000";
		ram_buffer(12054) := X"00000000";
		ram_buffer(12055) := X"00000000";
		ram_buffer(12056) := X"00000000";
		ram_buffer(12057) := X"00000000";
		ram_buffer(12058) := X"00000000";
		ram_buffer(12059) := X"00000000";
		ram_buffer(12060) := X"00000000";
		ram_buffer(12061) := X"00000000";
		ram_buffer(12062) := X"00000000";
		ram_buffer(12063) := X"00000000";
		ram_buffer(12064) := X"00000000";
		ram_buffer(12065) := X"00000000";
		ram_buffer(12066) := X"00000000";
		ram_buffer(12067) := X"00000000";
		ram_buffer(12068) := X"00000000";
		ram_buffer(12069) := X"00000000";
		ram_buffer(12070) := X"00000000";
		ram_buffer(12071) := X"00000000";
		ram_buffer(12072) := X"00000000";
		ram_buffer(12073) := X"00000000";
		ram_buffer(12074) := X"00000000";
		ram_buffer(12075) := X"00000000";
		ram_buffer(12076) := X"00000000";
		ram_buffer(12077) := X"00000000";
		ram_buffer(12078) := X"00000000";
		ram_buffer(12079) := X"00000000";
		ram_buffer(12080) := X"00000000";
		ram_buffer(12081) := X"00000000";
		ram_buffer(12082) := X"00000000";
		ram_buffer(12083) := X"00000000";
		ram_buffer(12084) := X"00000000";
		ram_buffer(12085) := X"00000000";
		ram_buffer(12086) := X"00000000";
		ram_buffer(12087) := X"00000000";
		ram_buffer(12088) := X"00000000";
		ram_buffer(12089) := X"00000000";
		ram_buffer(12090) := X"00000000";
		ram_buffer(12091) := X"00000000";
		ram_buffer(12092) := X"00000000";
		ram_buffer(12093) := X"00000000";
		ram_buffer(12094) := X"00000000";
		ram_buffer(12095) := X"00000000";
		ram_buffer(12096) := X"00000000";
		ram_buffer(12097) := X"00000000";
		ram_buffer(12098) := X"00000000";
		ram_buffer(12099) := X"00000000";
		ram_buffer(12100) := X"00000000";
		ram_buffer(12101) := X"00000000";
		ram_buffer(12102) := X"00000000";
		ram_buffer(12103) := X"00000000";
		ram_buffer(12104) := X"00000000";
		ram_buffer(12105) := X"00000000";
		ram_buffer(12106) := X"00000000";
		ram_buffer(12107) := X"00000000";
		ram_buffer(12108) := X"00000000";
		ram_buffer(12109) := X"00000000";
		ram_buffer(12110) := X"00000000";
		ram_buffer(12111) := X"00000000";
		ram_buffer(12112) := X"00000000";
		ram_buffer(12113) := X"00000000";
		ram_buffer(12114) := X"00000000";
		ram_buffer(12115) := X"00000000";
		ram_buffer(12116) := X"00000000";
		ram_buffer(12117) := X"00000000";
		ram_buffer(12118) := X"00000000";
		ram_buffer(12119) := X"00000000";
		ram_buffer(12120) := X"00000000";
		ram_buffer(12121) := X"00000000";
		ram_buffer(12122) := X"00000000";
		ram_buffer(12123) := X"00000000";
		ram_buffer(12124) := X"00000000";
		ram_buffer(12125) := X"00000000";
		ram_buffer(12126) := X"00000000";
		ram_buffer(12127) := X"00000000";
		ram_buffer(12128) := X"00000000";
		ram_buffer(12129) := X"00000000";
		ram_buffer(12130) := X"00000000";
		ram_buffer(12131) := X"00000000";
		ram_buffer(12132) := X"00000000";
		ram_buffer(12133) := X"00000000";
		ram_buffer(12134) := X"00000000";
		ram_buffer(12135) := X"00000000";
		ram_buffer(12136) := X"00000000";
		ram_buffer(12137) := X"00000000";
		ram_buffer(12138) := X"00000000";
		ram_buffer(12139) := X"00000000";
		ram_buffer(12140) := X"00000000";
		ram_buffer(12141) := X"00000000";
		ram_buffer(12142) := X"00000000";
		ram_buffer(12143) := X"00000000";
		ram_buffer(12144) := X"00000000";
		ram_buffer(12145) := X"00000000";
		ram_buffer(12146) := X"00000000";
		ram_buffer(12147) := X"00000000";
		ram_buffer(12148) := X"00000000";
		ram_buffer(12149) := X"00000000";
		ram_buffer(12150) := X"00000000";
		ram_buffer(12151) := X"00000000";
		ram_buffer(12152) := X"00000000";
		ram_buffer(12153) := X"00000000";
		ram_buffer(12154) := X"00000000";
		ram_buffer(12155) := X"00000000";
		ram_buffer(12156) := X"00000000";
		ram_buffer(12157) := X"00000000";
		ram_buffer(12158) := X"00000000";
		ram_buffer(12159) := X"00000000";
		ram_buffer(12160) := X"00000000";
		ram_buffer(12161) := X"00000000";
		ram_buffer(12162) := X"00000000";
		ram_buffer(12163) := X"00000000";
		ram_buffer(12164) := X"00000000";
		ram_buffer(12165) := X"00000000";
		ram_buffer(12166) := X"00000000";
		ram_buffer(12167) := X"00000000";
		ram_buffer(12168) := X"00000000";
		ram_buffer(12169) := X"00000000";
		ram_buffer(12170) := X"00000000";
		ram_buffer(12171) := X"00000000";
		ram_buffer(12172) := X"00000000";
		ram_buffer(12173) := X"00000000";
		ram_buffer(12174) := X"00000000";
		ram_buffer(12175) := X"00000000";
		ram_buffer(12176) := X"00000000";
		ram_buffer(12177) := X"00000000";
		ram_buffer(12178) := X"00000000";
		ram_buffer(12179) := X"00000000";
		ram_buffer(12180) := X"00000000";
		ram_buffer(12181) := X"00000000";
		ram_buffer(12182) := X"00000000";
		ram_buffer(12183) := X"00000000";
		ram_buffer(12184) := X"00000000";
		ram_buffer(12185) := X"00000000";
		ram_buffer(12186) := X"00000000";
		ram_buffer(12187) := X"00000000";
		ram_buffer(12188) := X"00000000";
		ram_buffer(12189) := X"00000000";
		ram_buffer(12190) := X"00000000";
		ram_buffer(12191) := X"00000000";
		ram_buffer(12192) := X"00000000";
		ram_buffer(12193) := X"00000000";
		ram_buffer(12194) := X"00000000";
		ram_buffer(12195) := X"00000000";
		ram_buffer(12196) := X"00000000";
		ram_buffer(12197) := X"00000000";
		ram_buffer(12198) := X"00000000";
		ram_buffer(12199) := X"00000000";
		ram_buffer(12200) := X"00000000";
		ram_buffer(12201) := X"00000000";
		ram_buffer(12202) := X"00000000";
		ram_buffer(12203) := X"00000000";
		ram_buffer(12204) := X"00000000";
		ram_buffer(12205) := X"00000000";
		ram_buffer(12206) := X"00000000";
		ram_buffer(12207) := X"00000000";
		ram_buffer(12208) := X"00000000";
		ram_buffer(12209) := X"00000000";
		ram_buffer(12210) := X"00000000";
		ram_buffer(12211) := X"00000000";
		ram_buffer(12212) := X"00000000";
		ram_buffer(12213) := X"00000000";
		ram_buffer(12214) := X"00000000";
		ram_buffer(12215) := X"00000000";
		ram_buffer(12216) := X"00000000";
		ram_buffer(12217) := X"00000000";
		ram_buffer(12218) := X"00000000";
		ram_buffer(12219) := X"00000000";
		ram_buffer(12220) := X"00000000";
		ram_buffer(12221) := X"00000000";
		ram_buffer(12222) := X"00000000";
		ram_buffer(12223) := X"00000000";
		ram_buffer(12224) := X"00000000";
		ram_buffer(12225) := X"00000000";
		ram_buffer(12226) := X"00000000";
		ram_buffer(12227) := X"00000000";
		ram_buffer(12228) := X"00000000";
		ram_buffer(12229) := X"00000000";
		ram_buffer(12230) := X"00000000";
		ram_buffer(12231) := X"00000000";
		ram_buffer(12232) := X"00000000";
		ram_buffer(12233) := X"00000000";
		ram_buffer(12234) := X"00000000";
		ram_buffer(12235) := X"00000000";
		ram_buffer(12236) := X"00000000";
		ram_buffer(12237) := X"00000000";
		ram_buffer(12238) := X"00000000";
		ram_buffer(12239) := X"00000000";
		ram_buffer(12240) := X"00000000";
		ram_buffer(12241) := X"00000000";
		ram_buffer(12242) := X"00000000";
		ram_buffer(12243) := X"00000000";
		ram_buffer(12244) := X"00000000";
		ram_buffer(12245) := X"00000000";
		ram_buffer(12246) := X"00000000";
		ram_buffer(12247) := X"00000000";
		ram_buffer(12248) := X"00000000";
		ram_buffer(12249) := X"00000000";
		ram_buffer(12250) := X"00000000";
		ram_buffer(12251) := X"00000000";
		ram_buffer(12252) := X"00000000";
		ram_buffer(12253) := X"00000000";
		ram_buffer(12254) := X"00000000";
		ram_buffer(12255) := X"00000000";
		ram_buffer(12256) := X"00000000";
		ram_buffer(12257) := X"00000000";
		ram_buffer(12258) := X"00000000";
		ram_buffer(12259) := X"00000000";
		ram_buffer(12260) := X"00000000";
		ram_buffer(12261) := X"00000000";
		ram_buffer(12262) := X"00000000";
		ram_buffer(12263) := X"00000000";
		ram_buffer(12264) := X"00000000";
		ram_buffer(12265) := X"00000000";
		ram_buffer(12266) := X"00000000";
		ram_buffer(12267) := X"00000000";
		ram_buffer(12268) := X"00000000";
		ram_buffer(12269) := X"00000000";
		ram_buffer(12270) := X"00000000";
		ram_buffer(12271) := X"00000000";
		ram_buffer(12272) := X"00000000";
		ram_buffer(12273) := X"00000000";
		ram_buffer(12274) := X"00000000";
		ram_buffer(12275) := X"00000000";
		ram_buffer(12276) := X"00000000";
		ram_buffer(12277) := X"00000000";
		ram_buffer(12278) := X"00000000";
		ram_buffer(12279) := X"00000000";
		ram_buffer(12280) := X"00000000";
		ram_buffer(12281) := X"00000000";
		ram_buffer(12282) := X"00000000";
		ram_buffer(12283) := X"00000000";
		ram_buffer(12284) := X"00000000";
		ram_buffer(12285) := X"00000000";
		ram_buffer(12286) := X"00000000";
		ram_buffer(12287) := X"00000000";
		ram_buffer(12288) := X"00000000";
		ram_buffer(12289) := X"00000000";
		ram_buffer(12290) := X"00000000";
		ram_buffer(12291) := X"00000000";
		ram_buffer(12292) := X"00000000";
		ram_buffer(12293) := X"00000000";
		ram_buffer(12294) := X"00000000";
		ram_buffer(12295) := X"00000000";
		ram_buffer(12296) := X"00000000";
		ram_buffer(12297) := X"00000000";
		ram_buffer(12298) := X"00000000";
		ram_buffer(12299) := X"00000000";
		ram_buffer(12300) := X"00000000";
		ram_buffer(12301) := X"00000000";
		ram_buffer(12302) := X"00000000";
		ram_buffer(12303) := X"00000000";
		ram_buffer(12304) := X"00000000";
		ram_buffer(12305) := X"00000000";
		ram_buffer(12306) := X"00000000";
		ram_buffer(12307) := X"00000000";
		ram_buffer(12308) := X"00000000";
		ram_buffer(12309) := X"00000000";
		ram_buffer(12310) := X"00000000";
		ram_buffer(12311) := X"00000000";
		ram_buffer(12312) := X"00000000";
		ram_buffer(12313) := X"00000000";
		ram_buffer(12314) := X"00000000";
		ram_buffer(12315) := X"00000000";
		ram_buffer(12316) := X"00000000";
		ram_buffer(12317) := X"00000000";
		ram_buffer(12318) := X"00000000";
		ram_buffer(12319) := X"00000000";
		ram_buffer(12320) := X"00000000";
		ram_buffer(12321) := X"00000000";
		ram_buffer(12322) := X"00000000";
		ram_buffer(12323) := X"00000000";
		ram_buffer(12324) := X"00000000";
		ram_buffer(12325) := X"00000000";
		ram_buffer(12326) := X"00000000";
		ram_buffer(12327) := X"00000000";
		ram_buffer(12328) := X"00000000";
		ram_buffer(12329) := X"00000000";
		ram_buffer(12330) := X"00000000";
		ram_buffer(12331) := X"00000000";
		ram_buffer(12332) := X"00000000";
		ram_buffer(12333) := X"00000000";
		ram_buffer(12334) := X"00000000";
		ram_buffer(12335) := X"00000000";
		ram_buffer(12336) := X"00000000";
		ram_buffer(12337) := X"00000000";
		ram_buffer(12338) := X"00000000";
		ram_buffer(12339) := X"00000000";
		ram_buffer(12340) := X"00000000";
		ram_buffer(12341) := X"00000000";
		ram_buffer(12342) := X"00000000";
		ram_buffer(12343) := X"00000000";
		ram_buffer(12344) := X"00000000";
		ram_buffer(12345) := X"00000000";
		ram_buffer(12346) := X"00000000";
		ram_buffer(12347) := X"00000000";
		ram_buffer(12348) := X"00000000";
		ram_buffer(12349) := X"00000000";
		ram_buffer(12350) := X"00000000";
		ram_buffer(12351) := X"00000000";
		ram_buffer(12352) := X"00000000";
		ram_buffer(12353) := X"00000000";
		ram_buffer(12354) := X"00000000";
		ram_buffer(12355) := X"00000000";
		ram_buffer(12356) := X"00000000";
		ram_buffer(12357) := X"00000000";
		ram_buffer(12358) := X"00000000";
		ram_buffer(12359) := X"00000000";
		ram_buffer(12360) := X"00000000";
		ram_buffer(12361) := X"00000000";
		ram_buffer(12362) := X"00000000";
		ram_buffer(12363) := X"00000000";
		ram_buffer(12364) := X"00000000";
		ram_buffer(12365) := X"00000000";
		ram_buffer(12366) := X"00000000";
		ram_buffer(12367) := X"00000000";
		ram_buffer(12368) := X"00000000";
		ram_buffer(12369) := X"00000000";
		ram_buffer(12370) := X"00000000";
		ram_buffer(12371) := X"00000000";
		ram_buffer(12372) := X"00000000";
		ram_buffer(12373) := X"00000000";
		ram_buffer(12374) := X"00000000";
		ram_buffer(12375) := X"00000000";
		ram_buffer(12376) := X"00000000";
		ram_buffer(12377) := X"00000000";
		ram_buffer(12378) := X"00000000";
		ram_buffer(12379) := X"00000000";
		ram_buffer(12380) := X"00000000";
		ram_buffer(12381) := X"00000000";
		ram_buffer(12382) := X"00000000";
		ram_buffer(12383) := X"00000000";
		ram_buffer(12384) := X"00000000";
		ram_buffer(12385) := X"00000000";
		ram_buffer(12386) := X"00000000";
		ram_buffer(12387) := X"00000000";
		ram_buffer(12388) := X"00000000";
		ram_buffer(12389) := X"00000000";
		ram_buffer(12390) := X"00000000";
		ram_buffer(12391) := X"00000000";
		ram_buffer(12392) := X"00000000";
		ram_buffer(12393) := X"00000000";
		ram_buffer(12394) := X"00000000";
		ram_buffer(12395) := X"00000000";
		ram_buffer(12396) := X"00000000";
		ram_buffer(12397) := X"00000000";
		ram_buffer(12398) := X"00000000";
		ram_buffer(12399) := X"00000000";
		ram_buffer(12400) := X"00000000";
		ram_buffer(12401) := X"00000000";
		ram_buffer(12402) := X"00000000";
		ram_buffer(12403) := X"00000000";
		ram_buffer(12404) := X"00000000";
		ram_buffer(12405) := X"00000000";
		ram_buffer(12406) := X"00000000";
		ram_buffer(12407) := X"00000000";
		ram_buffer(12408) := X"00000000";
		ram_buffer(12409) := X"00000000";
		ram_buffer(12410) := X"00000000";
		ram_buffer(12411) := X"00000000";
		ram_buffer(12412) := X"00000000";
		ram_buffer(12413) := X"00000000";
		ram_buffer(12414) := X"00000000";
		ram_buffer(12415) := X"00000000";
		ram_buffer(12416) := X"00000000";
		ram_buffer(12417) := X"00000000";
		ram_buffer(12418) := X"00000000";
		ram_buffer(12419) := X"00000000";
		ram_buffer(12420) := X"00000000";
		ram_buffer(12421) := X"00000000";
		ram_buffer(12422) := X"00000000";
		ram_buffer(12423) := X"00000000";
		ram_buffer(12424) := X"00000000";
		ram_buffer(12425) := X"00000000";
		ram_buffer(12426) := X"00000000";
		ram_buffer(12427) := X"00000000";
		ram_buffer(12428) := X"00000000";
		ram_buffer(12429) := X"00000000";
		ram_buffer(12430) := X"00000000";
		ram_buffer(12431) := X"00000000";
		ram_buffer(12432) := X"00000000";
		ram_buffer(12433) := X"00000000";
		ram_buffer(12434) := X"00000000";
		ram_buffer(12435) := X"00000000";
		ram_buffer(12436) := X"00000000";
		ram_buffer(12437) := X"00000000";
		ram_buffer(12438) := X"00000000";
		ram_buffer(12439) := X"00000000";
		ram_buffer(12440) := X"00000000";
		ram_buffer(12441) := X"00000000";
		ram_buffer(12442) := X"00000000";
		ram_buffer(12443) := X"00000000";
		ram_buffer(12444) := X"00000000";
		ram_buffer(12445) := X"00000000";
		ram_buffer(12446) := X"00000000";
		ram_buffer(12447) := X"00000000";
		ram_buffer(12448) := X"00000000";
		ram_buffer(12449) := X"00000000";
		ram_buffer(12450) := X"00000000";
		ram_buffer(12451) := X"00000000";
		ram_buffer(12452) := X"00000000";
		ram_buffer(12453) := X"00000000";
		ram_buffer(12454) := X"00000000";
		ram_buffer(12455) := X"00000000";
		ram_buffer(12456) := X"00000000";
		ram_buffer(12457) := X"00000000";
		ram_buffer(12458) := X"00000000";
		ram_buffer(12459) := X"00000000";
		ram_buffer(12460) := X"00000000";
		ram_buffer(12461) := X"00000000";
		ram_buffer(12462) := X"00000000";
		ram_buffer(12463) := X"00000000";
		ram_buffer(12464) := X"00000000";
		ram_buffer(12465) := X"00000000";
		ram_buffer(12466) := X"00000000";
		ram_buffer(12467) := X"00000000";
		ram_buffer(12468) := X"00000000";
		ram_buffer(12469) := X"00000000";
		ram_buffer(12470) := X"00000000";
		ram_buffer(12471) := X"00000000";
		ram_buffer(12472) := X"00000000";
		ram_buffer(12473) := X"00000000";
		ram_buffer(12474) := X"00000000";
		ram_buffer(12475) := X"00000000";
		ram_buffer(12476) := X"00000000";
		ram_buffer(12477) := X"00000000";
		ram_buffer(12478) := X"00000000";
		ram_buffer(12479) := X"00000000";
		ram_buffer(12480) := X"00000000";
		ram_buffer(12481) := X"00000000";
		ram_buffer(12482) := X"00000000";
		ram_buffer(12483) := X"00000000";
		ram_buffer(12484) := X"00000000";
		ram_buffer(12485) := X"00000000";
		ram_buffer(12486) := X"00000000";
		ram_buffer(12487) := X"00000000";
		ram_buffer(12488) := X"00000000";
		ram_buffer(12489) := X"00000000";
		ram_buffer(12490) := X"00000000";
		ram_buffer(12491) := X"00000000";
		ram_buffer(12492) := X"00000000";
		ram_buffer(12493) := X"00000000";
		ram_buffer(12494) := X"00000000";
		ram_buffer(12495) := X"00000000";
		ram_buffer(12496) := X"00000000";
		ram_buffer(12497) := X"00000000";
		ram_buffer(12498) := X"00000000";
		ram_buffer(12499) := X"00000000";
		ram_buffer(12500) := X"00000000";
		ram_buffer(12501) := X"00000000";
		ram_buffer(12502) := X"00000000";
		ram_buffer(12503) := X"00000000";
		ram_buffer(12504) := X"00000000";
		ram_buffer(12505) := X"00000000";
		ram_buffer(12506) := X"00000000";
		ram_buffer(12507) := X"00000000";
		ram_buffer(12508) := X"00000000";
		ram_buffer(12509) := X"00000000";
		ram_buffer(12510) := X"00000000";
		ram_buffer(12511) := X"00000000";
		ram_buffer(12512) := X"00000000";
		ram_buffer(12513) := X"00000000";
		ram_buffer(12514) := X"00000000";
		ram_buffer(12515) := X"00000000";
		ram_buffer(12516) := X"00000000";
		ram_buffer(12517) := X"00000000";
		ram_buffer(12518) := X"00000000";
		ram_buffer(12519) := X"00000000";
		ram_buffer(12520) := X"00000000";
		ram_buffer(12521) := X"00000000";
		ram_buffer(12522) := X"00000000";
		ram_buffer(12523) := X"00000000";
		ram_buffer(12524) := X"00000000";
		ram_buffer(12525) := X"00000000";
		ram_buffer(12526) := X"00000000";
		ram_buffer(12527) := X"00000000";
		ram_buffer(12528) := X"00000000";
		ram_buffer(12529) := X"00000000";
		ram_buffer(12530) := X"00000000";
		ram_buffer(12531) := X"00000000";
		ram_buffer(12532) := X"00000000";
		ram_buffer(12533) := X"00000000";
		ram_buffer(12534) := X"00000000";
		ram_buffer(12535) := X"00000000";
		ram_buffer(12536) := X"00000000";
		ram_buffer(12537) := X"00000000";
		ram_buffer(12538) := X"00000000";
		ram_buffer(12539) := X"00000000";
		ram_buffer(12540) := X"00000000";
		ram_buffer(12541) := X"00000000";
		ram_buffer(12542) := X"00000000";
		ram_buffer(12543) := X"00000000";
		ram_buffer(12544) := X"00000000";
		ram_buffer(12545) := X"00000000";
		ram_buffer(12546) := X"00000000";
		ram_buffer(12547) := X"00000000";
		ram_buffer(12548) := X"00000000";
		ram_buffer(12549) := X"00000000";
		ram_buffer(12550) := X"00000000";
		ram_buffer(12551) := X"00000000";
		ram_buffer(12552) := X"00000000";
		ram_buffer(12553) := X"00000000";
		ram_buffer(12554) := X"00000000";
		ram_buffer(12555) := X"00000000";
		ram_buffer(12556) := X"00000000";
		ram_buffer(12557) := X"00000000";
		ram_buffer(12558) := X"00000000";
		ram_buffer(12559) := X"00000000";
		ram_buffer(12560) := X"00000000";
		ram_buffer(12561) := X"00000000";
		ram_buffer(12562) := X"00000000";
		ram_buffer(12563) := X"00000000";
		ram_buffer(12564) := X"00000000";
		ram_buffer(12565) := X"00000000";
		ram_buffer(12566) := X"00000000";
		ram_buffer(12567) := X"00000000";
		ram_buffer(12568) := X"00000000";
		ram_buffer(12569) := X"00000000";
		ram_buffer(12570) := X"00000000";
		ram_buffer(12571) := X"00000000";
		ram_buffer(12572) := X"00000000";
		ram_buffer(12573) := X"00000000";
		ram_buffer(12574) := X"00000000";
		ram_buffer(12575) := X"00000000";
		ram_buffer(12576) := X"00000000";
		ram_buffer(12577) := X"00000000";
		ram_buffer(12578) := X"00000000";
		ram_buffer(12579) := X"00000000";
		ram_buffer(12580) := X"00000000";
		ram_buffer(12581) := X"00000000";
		ram_buffer(12582) := X"00000000";
		ram_buffer(12583) := X"00000000";
		ram_buffer(12584) := X"00000000";
		ram_buffer(12585) := X"00000000";
		ram_buffer(12586) := X"00000000";
		ram_buffer(12587) := X"00000000";
		ram_buffer(12588) := X"00000000";
		ram_buffer(12589) := X"00000000";
		ram_buffer(12590) := X"00000000";
		ram_buffer(12591) := X"00000000";
		ram_buffer(12592) := X"00000000";
		ram_buffer(12593) := X"00000000";
		ram_buffer(12594) := X"00000000";
		ram_buffer(12595) := X"00000000";
		ram_buffer(12596) := X"00000000";
		ram_buffer(12597) := X"00000000";
		ram_buffer(12598) := X"00000000";
		ram_buffer(12599) := X"00000000";
		ram_buffer(12600) := X"00000000";
		ram_buffer(12601) := X"00000000";
		ram_buffer(12602) := X"00000000";
		ram_buffer(12603) := X"00000000";
		ram_buffer(12604) := X"00000000";
		ram_buffer(12605) := X"00000000";
		ram_buffer(12606) := X"00000000";
		ram_buffer(12607) := X"00000000";
		ram_buffer(12608) := X"00000000";
		ram_buffer(12609) := X"00000000";
		ram_buffer(12610) := X"00000000";
		ram_buffer(12611) := X"00000000";
		ram_buffer(12612) := X"00000000";
		ram_buffer(12613) := X"00000000";
		ram_buffer(12614) := X"00000000";
		ram_buffer(12615) := X"00000000";
		ram_buffer(12616) := X"00000000";
		ram_buffer(12617) := X"00000000";
		ram_buffer(12618) := X"00000000";
		ram_buffer(12619) := X"00000000";
		ram_buffer(12620) := X"00000000";
		ram_buffer(12621) := X"00000000";
		ram_buffer(12622) := X"00000000";
		ram_buffer(12623) := X"00000000";
		ram_buffer(12624) := X"00000000";
		ram_buffer(12625) := X"00000000";
		ram_buffer(12626) := X"00000000";
		ram_buffer(12627) := X"00000000";
		ram_buffer(12628) := X"00000000";
		ram_buffer(12629) := X"00000000";
		ram_buffer(12630) := X"00000000";
		ram_buffer(12631) := X"00000000";
		ram_buffer(12632) := X"00000000";
		ram_buffer(12633) := X"00000000";
		ram_buffer(12634) := X"00000000";
		ram_buffer(12635) := X"00000000";
		ram_buffer(12636) := X"00000000";
		ram_buffer(12637) := X"00000000";
		ram_buffer(12638) := X"00000000";
		ram_buffer(12639) := X"00000000";
		ram_buffer(12640) := X"00000000";
		ram_buffer(12641) := X"00000000";
		ram_buffer(12642) := X"00000000";
		ram_buffer(12643) := X"00000000";
		ram_buffer(12644) := X"00000000";
		ram_buffer(12645) := X"00000000";
		ram_buffer(12646) := X"00000000";
		ram_buffer(12647) := X"00000000";
		ram_buffer(12648) := X"00000000";
		ram_buffer(12649) := X"00000000";
		ram_buffer(12650) := X"00000000";
		ram_buffer(12651) := X"00000000";
		ram_buffer(12652) := X"00000000";
		ram_buffer(12653) := X"00000000";
		ram_buffer(12654) := X"00000000";
		ram_buffer(12655) := X"00000000";
		ram_buffer(12656) := X"00000000";
		ram_buffer(12657) := X"00000000";
		ram_buffer(12658) := X"00000000";
		ram_buffer(12659) := X"00000000";
		ram_buffer(12660) := X"00000000";
		ram_buffer(12661) := X"00000000";
		ram_buffer(12662) := X"00000000";
		ram_buffer(12663) := X"00000000";
		ram_buffer(12664) := X"00000000";
		ram_buffer(12665) := X"00000000";
		ram_buffer(12666) := X"00000000";
		ram_buffer(12667) := X"00000000";
		ram_buffer(12668) := X"00000000";
		ram_buffer(12669) := X"00000000";
		ram_buffer(12670) := X"00000000";
		ram_buffer(12671) := X"00000000";
		ram_buffer(12672) := X"00000000";
		ram_buffer(12673) := X"00000000";
		ram_buffer(12674) := X"00000000";
		ram_buffer(12675) := X"00000000";
		ram_buffer(12676) := X"00000000";
		ram_buffer(12677) := X"00000000";
		ram_buffer(12678) := X"00000000";
		ram_buffer(12679) := X"00000000";
		ram_buffer(12680) := X"00000000";
		ram_buffer(12681) := X"00000000";
		ram_buffer(12682) := X"00000000";
		ram_buffer(12683) := X"00000000";
		ram_buffer(12684) := X"00000000";
		ram_buffer(12685) := X"00000000";
		ram_buffer(12686) := X"00000000";
		ram_buffer(12687) := X"00000000";
		ram_buffer(12688) := X"00000000";
		ram_buffer(12689) := X"00000000";
		ram_buffer(12690) := X"00000000";
		ram_buffer(12691) := X"00000000";
		ram_buffer(12692) := X"00000000";
		ram_buffer(12693) := X"00000000";
		ram_buffer(12694) := X"00000000";
		ram_buffer(12695) := X"00000000";
		ram_buffer(12696) := X"00000000";
		ram_buffer(12697) := X"00000000";
		ram_buffer(12698) := X"00000000";
		ram_buffer(12699) := X"00000000";
		ram_buffer(12700) := X"00000000";
		ram_buffer(12701) := X"00000000";
		ram_buffer(12702) := X"00000000";
		ram_buffer(12703) := X"00000000";
		ram_buffer(12704) := X"00000000";
		ram_buffer(12705) := X"00000000";
		ram_buffer(12706) := X"00000000";
		ram_buffer(12707) := X"00000000";
		ram_buffer(12708) := X"00000000";
		ram_buffer(12709) := X"00000000";
		ram_buffer(12710) := X"00000000";
		ram_buffer(12711) := X"00000000";
		ram_buffer(12712) := X"00000000";
		ram_buffer(12713) := X"00000000";
		ram_buffer(12714) := X"00000000";
		ram_buffer(12715) := X"00000000";
		ram_buffer(12716) := X"00000000";
		ram_buffer(12717) := X"00000000";
		ram_buffer(12718) := X"00000000";
		ram_buffer(12719) := X"00000000";
		ram_buffer(12720) := X"00000000";
		ram_buffer(12721) := X"00000000";
		ram_buffer(12722) := X"00000000";
		ram_buffer(12723) := X"00000000";
		ram_buffer(12724) := X"00000000";
		ram_buffer(12725) := X"00000000";
		ram_buffer(12726) := X"00000000";
		ram_buffer(12727) := X"00000000";
		ram_buffer(12728) := X"00000000";
		ram_buffer(12729) := X"00000000";
		ram_buffer(12730) := X"00000000";
		ram_buffer(12731) := X"00000000";
		ram_buffer(12732) := X"00000000";
		ram_buffer(12733) := X"00000000";
		ram_buffer(12734) := X"00000000";
		ram_buffer(12735) := X"00000000";
		ram_buffer(12736) := X"00000000";
		ram_buffer(12737) := X"00000000";
		ram_buffer(12738) := X"00000000";
		ram_buffer(12739) := X"00000000";
		ram_buffer(12740) := X"00000000";
		ram_buffer(12741) := X"00000000";
		ram_buffer(12742) := X"00000000";
		ram_buffer(12743) := X"00000000";
		ram_buffer(12744) := X"00000000";
		ram_buffer(12745) := X"00000000";
		ram_buffer(12746) := X"00000000";
		ram_buffer(12747) := X"00000000";
		ram_buffer(12748) := X"00000000";
		ram_buffer(12749) := X"00000000";
		ram_buffer(12750) := X"00000000";
		ram_buffer(12751) := X"00000000";
		ram_buffer(12752) := X"00000000";
		ram_buffer(12753) := X"00000000";
		ram_buffer(12754) := X"00000000";
		ram_buffer(12755) := X"00000000";
		ram_buffer(12756) := X"00000000";
		ram_buffer(12757) := X"00000000";
		ram_buffer(12758) := X"00000000";
		ram_buffer(12759) := X"00000000";
		ram_buffer(12760) := X"00000000";
		ram_buffer(12761) := X"00000000";
		ram_buffer(12762) := X"00000000";
		ram_buffer(12763) := X"00000000";
		ram_buffer(12764) := X"00000000";
		ram_buffer(12765) := X"00000000";
		ram_buffer(12766) := X"00000000";
		ram_buffer(12767) := X"00000000";
		ram_buffer(12768) := X"00000000";
		ram_buffer(12769) := X"00000000";
		ram_buffer(12770) := X"00000000";
		ram_buffer(12771) := X"00000000";
		ram_buffer(12772) := X"00000000";
		ram_buffer(12773) := X"00000000";
		ram_buffer(12774) := X"00000000";
		ram_buffer(12775) := X"00000000";
		ram_buffer(12776) := X"00000000";
		ram_buffer(12777) := X"00000000";
		ram_buffer(12778) := X"00000000";
		ram_buffer(12779) := X"00000000";
		ram_buffer(12780) := X"00000000";
		ram_buffer(12781) := X"00000000";
		ram_buffer(12782) := X"00000000";
		ram_buffer(12783) := X"00000000";
		ram_buffer(12784) := X"00000000";
		ram_buffer(12785) := X"00000000";
		ram_buffer(12786) := X"00000000";
		ram_buffer(12787) := X"00000000";
		ram_buffer(12788) := X"00000000";
		ram_buffer(12789) := X"00000000";
		ram_buffer(12790) := X"00000000";
		ram_buffer(12791) := X"00000000";
		ram_buffer(12792) := X"00000000";
		ram_buffer(12793) := X"00000000";
		ram_buffer(12794) := X"00000000";
		ram_buffer(12795) := X"00000000";
		ram_buffer(12796) := X"00000000";
		ram_buffer(12797) := X"00000000";
		ram_buffer(12798) := X"00000000";
		ram_buffer(12799) := X"00000000";
		ram_buffer(12800) := X"00000000";
		ram_buffer(12801) := X"00000000";
		ram_buffer(12802) := X"00000000";
		ram_buffer(12803) := X"00000000";
		ram_buffer(12804) := X"00000000";
		ram_buffer(12805) := X"00000000";
		ram_buffer(12806) := X"00000000";
		ram_buffer(12807) := X"00000000";
		ram_buffer(12808) := X"00000000";
		ram_buffer(12809) := X"00000000";
		ram_buffer(12810) := X"00000000";
		ram_buffer(12811) := X"00000000";
		ram_buffer(12812) := X"00000000";
		ram_buffer(12813) := X"00000000";
		ram_buffer(12814) := X"00000000";
		ram_buffer(12815) := X"00000000";
		ram_buffer(12816) := X"00000000";
		ram_buffer(12817) := X"00000000";
		ram_buffer(12818) := X"00000000";
		ram_buffer(12819) := X"00000000";
		ram_buffer(12820) := X"00000000";
		ram_buffer(12821) := X"00000000";
		ram_buffer(12822) := X"00000000";
		ram_buffer(12823) := X"00000000";
		ram_buffer(12824) := X"00000000";
		ram_buffer(12825) := X"00000000";
		ram_buffer(12826) := X"00000000";
		ram_buffer(12827) := X"00000000";
		ram_buffer(12828) := X"00000000";
		ram_buffer(12829) := X"00000000";
		ram_buffer(12830) := X"00000000";
		ram_buffer(12831) := X"00000000";
		ram_buffer(12832) := X"00000000";
		ram_buffer(12833) := X"00000000";
		ram_buffer(12834) := X"00000000";
		ram_buffer(12835) := X"00000000";
		ram_buffer(12836) := X"00000000";
		ram_buffer(12837) := X"00000000";
		ram_buffer(12838) := X"00000000";
		ram_buffer(12839) := X"00000000";
		ram_buffer(12840) := X"00000000";
		ram_buffer(12841) := X"00000000";
		ram_buffer(12842) := X"00000000";
		ram_buffer(12843) := X"00000000";
		ram_buffer(12844) := X"00000000";
		ram_buffer(12845) := X"00000000";
		ram_buffer(12846) := X"00000000";
		ram_buffer(12847) := X"00000000";
		ram_buffer(12848) := X"00000000";
		ram_buffer(12849) := X"00000000";
		ram_buffer(12850) := X"00000000";
		ram_buffer(12851) := X"00000000";
		ram_buffer(12852) := X"00000000";
		ram_buffer(12853) := X"00000000";
		ram_buffer(12854) := X"00000000";
		ram_buffer(12855) := X"00000000";
		ram_buffer(12856) := X"00000000";
		ram_buffer(12857) := X"00000000";
		ram_buffer(12858) := X"00000000";
		ram_buffer(12859) := X"00000000";
		ram_buffer(12860) := X"00000000";
		ram_buffer(12861) := X"00000000";
		ram_buffer(12862) := X"00000000";
		ram_buffer(12863) := X"00000000";
		ram_buffer(12864) := X"00000000";
		ram_buffer(12865) := X"00000000";
		ram_buffer(12866) := X"00000000";
		ram_buffer(12867) := X"00000000";
		ram_buffer(12868) := X"00000000";
		ram_buffer(12869) := X"00000000";
		ram_buffer(12870) := X"00000000";
		ram_buffer(12871) := X"00000000";
		ram_buffer(12872) := X"00000000";
		ram_buffer(12873) := X"00000000";
		ram_buffer(12874) := X"00000000";
		ram_buffer(12875) := X"00000000";
		ram_buffer(12876) := X"00000000";
		ram_buffer(12877) := X"00000000";
		ram_buffer(12878) := X"00000000";
		ram_buffer(12879) := X"00000000";
		ram_buffer(12880) := X"00000000";
		ram_buffer(12881) := X"00000000";
		ram_buffer(12882) := X"00000000";
		ram_buffer(12883) := X"00000000";
		ram_buffer(12884) := X"00000000";
		ram_buffer(12885) := X"00000000";
		ram_buffer(12886) := X"00000000";
		ram_buffer(12887) := X"00000000";
		ram_buffer(12888) := X"00000000";
		ram_buffer(12889) := X"00000000";
		ram_buffer(12890) := X"00000000";
		ram_buffer(12891) := X"00000000";
		ram_buffer(12892) := X"00000000";
		ram_buffer(12893) := X"00000000";
		ram_buffer(12894) := X"00000000";
		ram_buffer(12895) := X"00000000";
		ram_buffer(12896) := X"00000000";
		ram_buffer(12897) := X"00000000";
		ram_buffer(12898) := X"00000000";
		ram_buffer(12899) := X"00000000";
		ram_buffer(12900) := X"00000000";
		ram_buffer(12901) := X"00000000";
		ram_buffer(12902) := X"00000000";
		ram_buffer(12903) := X"00000000";
		ram_buffer(12904) := X"00000000";
		ram_buffer(12905) := X"00000000";
		ram_buffer(12906) := X"00000000";
		ram_buffer(12907) := X"00000000";
		ram_buffer(12908) := X"00000000";
		ram_buffer(12909) := X"00000000";
		ram_buffer(12910) := X"00000000";
		ram_buffer(12911) := X"00000000";
		ram_buffer(12912) := X"00000000";
		ram_buffer(12913) := X"00000000";
		ram_buffer(12914) := X"00000000";
		ram_buffer(12915) := X"00000000";
		ram_buffer(12916) := X"00000000";
		ram_buffer(12917) := X"00000000";
		ram_buffer(12918) := X"00000000";
		ram_buffer(12919) := X"00000000";
		ram_buffer(12920) := X"00000000";
		ram_buffer(12921) := X"00000000";
		ram_buffer(12922) := X"00000000";
		ram_buffer(12923) := X"00000000";
		ram_buffer(12924) := X"00000000";
		ram_buffer(12925) := X"00000000";
		ram_buffer(12926) := X"00000000";
		ram_buffer(12927) := X"00000000";
		ram_buffer(12928) := X"00000000";
		ram_buffer(12929) := X"00000000";
		ram_buffer(12930) := X"00000000";
		ram_buffer(12931) := X"00000000";
		ram_buffer(12932) := X"00000000";
		ram_buffer(12933) := X"00000000";
		ram_buffer(12934) := X"00000000";
		ram_buffer(12935) := X"00000000";
		ram_buffer(12936) := X"00000000";
		ram_buffer(12937) := X"00000000";
		ram_buffer(12938) := X"00000000";
		ram_buffer(12939) := X"00000000";
		ram_buffer(12940) := X"00000000";
		ram_buffer(12941) := X"00000000";
		ram_buffer(12942) := X"00000000";
		ram_buffer(12943) := X"00000000";
		ram_buffer(12944) := X"00000000";
		ram_buffer(12945) := X"00000000";
		ram_buffer(12946) := X"00000000";
		ram_buffer(12947) := X"00000000";
		ram_buffer(12948) := X"00000000";
		ram_buffer(12949) := X"00000000";
		ram_buffer(12950) := X"00000000";
		ram_buffer(12951) := X"00000000";
		ram_buffer(12952) := X"00000000";
		ram_buffer(12953) := X"00000000";
		ram_buffer(12954) := X"00000000";
		ram_buffer(12955) := X"00000000";
		ram_buffer(12956) := X"00000000";
		ram_buffer(12957) := X"00000000";
		ram_buffer(12958) := X"00000000";
		ram_buffer(12959) := X"00000000";
		ram_buffer(12960) := X"00000000";
		ram_buffer(12961) := X"00000000";
		ram_buffer(12962) := X"00000000";
		ram_buffer(12963) := X"00000000";
		ram_buffer(12964) := X"00000000";
		ram_buffer(12965) := X"00000000";
		ram_buffer(12966) := X"00000000";
		ram_buffer(12967) := X"00000000";
		ram_buffer(12968) := X"00000000";
		ram_buffer(12969) := X"00000000";
		ram_buffer(12970) := X"00000000";
		ram_buffer(12971) := X"00000000";
		ram_buffer(12972) := X"00000000";
		ram_buffer(12973) := X"00000000";
		ram_buffer(12974) := X"00000000";
		ram_buffer(12975) := X"00000000";
		ram_buffer(12976) := X"00000000";
		ram_buffer(12977) := X"00000000";
		ram_buffer(12978) := X"00000000";
		ram_buffer(12979) := X"00000000";
		ram_buffer(12980) := X"00000000";
		ram_buffer(12981) := X"00000000";
		ram_buffer(12982) := X"00000000";
		ram_buffer(12983) := X"00000000";
		ram_buffer(12984) := X"00000000";
		ram_buffer(12985) := X"00000000";
		ram_buffer(12986) := X"00000000";
		ram_buffer(12987) := X"00000000";
		ram_buffer(12988) := X"00000000";
		ram_buffer(12989) := X"00000000";
		ram_buffer(12990) := X"00000000";
		ram_buffer(12991) := X"00000000";
		ram_buffer(12992) := X"00000000";
		ram_buffer(12993) := X"00000000";
		ram_buffer(12994) := X"00000000";
		ram_buffer(12995) := X"00000000";
		ram_buffer(12996) := X"00000000";
		ram_buffer(12997) := X"00000000";
		ram_buffer(12998) := X"00000000";
		ram_buffer(12999) := X"00000000";
		ram_buffer(13000) := X"00000000";
		ram_buffer(13001) := X"00000000";
		ram_buffer(13002) := X"00000000";
		ram_buffer(13003) := X"00000000";
		ram_buffer(13004) := X"00000000";
		ram_buffer(13005) := X"00000000";
		ram_buffer(13006) := X"00000000";
		ram_buffer(13007) := X"00000000";
		ram_buffer(13008) := X"00000000";
		ram_buffer(13009) := X"00000000";
		ram_buffer(13010) := X"00000000";
		ram_buffer(13011) := X"00000000";
		ram_buffer(13012) := X"00000000";
		ram_buffer(13013) := X"00000000";
		ram_buffer(13014) := X"00000000";
		ram_buffer(13015) := X"00000000";
		ram_buffer(13016) := X"00000000";
		ram_buffer(13017) := X"00000000";
		ram_buffer(13018) := X"00000000";
		ram_buffer(13019) := X"00000000";
		ram_buffer(13020) := X"00000000";
		ram_buffer(13021) := X"00000000";
		ram_buffer(13022) := X"00000000";
		ram_buffer(13023) := X"00000000";
		ram_buffer(13024) := X"00000000";
		ram_buffer(13025) := X"00000000";
		ram_buffer(13026) := X"00000000";
		ram_buffer(13027) := X"00000000";
		ram_buffer(13028) := X"00000000";
		ram_buffer(13029) := X"00000000";
		ram_buffer(13030) := X"00000000";
		ram_buffer(13031) := X"00000000";
		ram_buffer(13032) := X"00000000";
		ram_buffer(13033) := X"00000000";
		ram_buffer(13034) := X"00000000";
		ram_buffer(13035) := X"00000000";
		ram_buffer(13036) := X"00000000";
		ram_buffer(13037) := X"00000000";
		ram_buffer(13038) := X"00000000";
		ram_buffer(13039) := X"00000000";
		ram_buffer(13040) := X"00000000";
		ram_buffer(13041) := X"00000000";
		ram_buffer(13042) := X"00000000";
		ram_buffer(13043) := X"00000000";
		ram_buffer(13044) := X"00000000";
		ram_buffer(13045) := X"00000000";
		ram_buffer(13046) := X"00000000";
		ram_buffer(13047) := X"00000000";
		ram_buffer(13048) := X"00000000";
		ram_buffer(13049) := X"00000000";
		ram_buffer(13050) := X"00000000";
		ram_buffer(13051) := X"00000000";
		ram_buffer(13052) := X"00000000";
		ram_buffer(13053) := X"00000000";
		ram_buffer(13054) := X"00000000";
		ram_buffer(13055) := X"00000000";
		ram_buffer(13056) := X"00000000";
		ram_buffer(13057) := X"00000000";
		ram_buffer(13058) := X"00000000";
		ram_buffer(13059) := X"00000000";
		ram_buffer(13060) := X"00000000";
		ram_buffer(13061) := X"00000000";
		ram_buffer(13062) := X"00000000";
		ram_buffer(13063) := X"00000000";
		ram_buffer(13064) := X"00000000";
		ram_buffer(13065) := X"00000000";
		ram_buffer(13066) := X"00000000";
		ram_buffer(13067) := X"00000000";
		ram_buffer(13068) := X"00000000";
		ram_buffer(13069) := X"00000000";
		ram_buffer(13070) := X"00000000";
		ram_buffer(13071) := X"00000000";
		ram_buffer(13072) := X"00000000";
		ram_buffer(13073) := X"00000000";
		ram_buffer(13074) := X"00000000";
		ram_buffer(13075) := X"00000000";
		ram_buffer(13076) := X"00000000";
		ram_buffer(13077) := X"00000000";
		ram_buffer(13078) := X"00000000";
		ram_buffer(13079) := X"00000000";
		ram_buffer(13080) := X"00000000";
		ram_buffer(13081) := X"00000000";
		ram_buffer(13082) := X"00000000";
		ram_buffer(13083) := X"00000000";
		ram_buffer(13084) := X"00000000";
		ram_buffer(13085) := X"00000000";
		ram_buffer(13086) := X"00000000";
		ram_buffer(13087) := X"00000000";
		ram_buffer(13088) := X"00000000";
		ram_buffer(13089) := X"00000000";
		ram_buffer(13090) := X"00000000";
		ram_buffer(13091) := X"00000000";
		ram_buffer(13092) := X"00000000";
		ram_buffer(13093) := X"00000000";
		ram_buffer(13094) := X"00000000";
		ram_buffer(13095) := X"00000000";
		ram_buffer(13096) := X"00000000";
		ram_buffer(13097) := X"00000000";
		ram_buffer(13098) := X"00000000";
		ram_buffer(13099) := X"00000000";
		ram_buffer(13100) := X"00000000";
		ram_buffer(13101) := X"00000000";
		ram_buffer(13102) := X"00000000";
		ram_buffer(13103) := X"00000000";
		ram_buffer(13104) := X"00000000";
		ram_buffer(13105) := X"00000000";
		ram_buffer(13106) := X"00000000";
		ram_buffer(13107) := X"00000000";
		ram_buffer(13108) := X"00000000";
		ram_buffer(13109) := X"00000000";
		ram_buffer(13110) := X"00000000";
		ram_buffer(13111) := X"00000000";
		ram_buffer(13112) := X"00000000";
		ram_buffer(13113) := X"00000000";
		ram_buffer(13114) := X"00000000";
		ram_buffer(13115) := X"00000000";
		ram_buffer(13116) := X"00000000";
		ram_buffer(13117) := X"00000000";
		ram_buffer(13118) := X"00000000";
		ram_buffer(13119) := X"00000000";
		ram_buffer(13120) := X"00000000";
		ram_buffer(13121) := X"00000000";
		ram_buffer(13122) := X"00000000";
		ram_buffer(13123) := X"00000000";
		ram_buffer(13124) := X"00000000";
		ram_buffer(13125) := X"00000000";
		ram_buffer(13126) := X"00000000";
		ram_buffer(13127) := X"00000000";
		ram_buffer(13128) := X"00000000";
		ram_buffer(13129) := X"00000000";
		ram_buffer(13130) := X"00000000";
		ram_buffer(13131) := X"00000000";
		ram_buffer(13132) := X"00000000";
		ram_buffer(13133) := X"00000000";
		ram_buffer(13134) := X"00000000";
		ram_buffer(13135) := X"00000000";
		ram_buffer(13136) := X"00000000";
		ram_buffer(13137) := X"00000000";
		ram_buffer(13138) := X"00000000";
		ram_buffer(13139) := X"00000000";
		ram_buffer(13140) := X"00000000";
		ram_buffer(13141) := X"00000000";
		ram_buffer(13142) := X"00000000";
		ram_buffer(13143) := X"00000000";
		ram_buffer(13144) := X"00000000";
		ram_buffer(13145) := X"00000000";
		ram_buffer(13146) := X"00000000";
		ram_buffer(13147) := X"00000000";
		ram_buffer(13148) := X"00000000";
		ram_buffer(13149) := X"00000000";
		ram_buffer(13150) := X"00000000";
		ram_buffer(13151) := X"00000000";
		ram_buffer(13152) := X"00000000";
		ram_buffer(13153) := X"00000000";
		ram_buffer(13154) := X"00000000";
		ram_buffer(13155) := X"00000000";
		ram_buffer(13156) := X"00000000";
		ram_buffer(13157) := X"00000000";
		ram_buffer(13158) := X"00000000";
		ram_buffer(13159) := X"00000000";
		ram_buffer(13160) := X"00000000";
		ram_buffer(13161) := X"00000000";
		ram_buffer(13162) := X"00000000";
		ram_buffer(13163) := X"00000000";
		ram_buffer(13164) := X"00000000";
		ram_buffer(13165) := X"00000000";
		ram_buffer(13166) := X"00000000";
		ram_buffer(13167) := X"00000000";
		ram_buffer(13168) := X"00000000";
		ram_buffer(13169) := X"00000000";
		ram_buffer(13170) := X"00000000";
		ram_buffer(13171) := X"00000000";
		ram_buffer(13172) := X"00000000";
		ram_buffer(13173) := X"00000000";
		ram_buffer(13174) := X"00000000";
		ram_buffer(13175) := X"00000000";
		ram_buffer(13176) := X"00000000";
		ram_buffer(13177) := X"00000000";
		ram_buffer(13178) := X"00000000";
		ram_buffer(13179) := X"00000000";
		ram_buffer(13180) := X"00000000";
		ram_buffer(13181) := X"00000000";
		ram_buffer(13182) := X"00000000";
		ram_buffer(13183) := X"00000000";
		ram_buffer(13184) := X"00000000";
		ram_buffer(13185) := X"00000000";
		ram_buffer(13186) := X"00000000";
		ram_buffer(13187) := X"00000000";
		ram_buffer(13188) := X"00000000";
		ram_buffer(13189) := X"00000000";
		ram_buffer(13190) := X"00000000";
		ram_buffer(13191) := X"00000000";
		ram_buffer(13192) := X"00000000";
		ram_buffer(13193) := X"00000000";
		ram_buffer(13194) := X"00000000";
		ram_buffer(13195) := X"00000000";
		ram_buffer(13196) := X"00000000";
		ram_buffer(13197) := X"00000000";
		ram_buffer(13198) := X"00000000";
		ram_buffer(13199) := X"00000000";
		ram_buffer(13200) := X"00000000";
		ram_buffer(13201) := X"00000000";
		ram_buffer(13202) := X"00000000";
		ram_buffer(13203) := X"00000000";
		ram_buffer(13204) := X"00000000";
		ram_buffer(13205) := X"00000000";
		ram_buffer(13206) := X"00000000";
		ram_buffer(13207) := X"00000000";
		ram_buffer(13208) := X"00000000";
		ram_buffer(13209) := X"00000000";
		ram_buffer(13210) := X"00000000";
		ram_buffer(13211) := X"00000000";
		ram_buffer(13212) := X"00000000";
		ram_buffer(13213) := X"00000000";
		ram_buffer(13214) := X"00000000";
		ram_buffer(13215) := X"00000000";
		ram_buffer(13216) := X"00000000";
		ram_buffer(13217) := X"00000000";
		ram_buffer(13218) := X"00000000";
		ram_buffer(13219) := X"00000000";
		ram_buffer(13220) := X"00000000";
		ram_buffer(13221) := X"00000000";
		ram_buffer(13222) := X"00000000";
		ram_buffer(13223) := X"00000000";
		ram_buffer(13224) := X"00000000";
		ram_buffer(13225) := X"00000000";
		ram_buffer(13226) := X"00000000";
		ram_buffer(13227) := X"00000000";
		ram_buffer(13228) := X"00000000";
		ram_buffer(13229) := X"00000000";
		ram_buffer(13230) := X"00000000";
		ram_buffer(13231) := X"00000000";
		ram_buffer(13232) := X"00000000";
		ram_buffer(13233) := X"00000000";
		ram_buffer(13234) := X"00000000";
		ram_buffer(13235) := X"00000000";
		ram_buffer(13236) := X"00000000";
		ram_buffer(13237) := X"00000000";
		ram_buffer(13238) := X"00000000";
		ram_buffer(13239) := X"00000000";
		ram_buffer(13240) := X"00000000";
		ram_buffer(13241) := X"00000000";
		ram_buffer(13242) := X"00000000";
		ram_buffer(13243) := X"00000000";
		ram_buffer(13244) := X"00000000";
		ram_buffer(13245) := X"00000000";
		ram_buffer(13246) := X"00000000";
		ram_buffer(13247) := X"00000000";
		ram_buffer(13248) := X"00000000";
		ram_buffer(13249) := X"00000000";
		ram_buffer(13250) := X"00000000";
		ram_buffer(13251) := X"00000000";
		ram_buffer(13252) := X"00000000";
		ram_buffer(13253) := X"00000000";
		ram_buffer(13254) := X"00000000";
		ram_buffer(13255) := X"00000000";
		ram_buffer(13256) := X"00000000";
		ram_buffer(13257) := X"00000000";
		ram_buffer(13258) := X"00000000";
		ram_buffer(13259) := X"00000000";
		ram_buffer(13260) := X"00000000";
		ram_buffer(13261) := X"00000000";
		ram_buffer(13262) := X"00000000";
		ram_buffer(13263) := X"00000000";
		ram_buffer(13264) := X"00000000";
		ram_buffer(13265) := X"00000000";
		ram_buffer(13266) := X"00000000";
		ram_buffer(13267) := X"00000000";
		ram_buffer(13268) := X"00000000";
		ram_buffer(13269) := X"00000000";
		ram_buffer(13270) := X"00000000";
		ram_buffer(13271) := X"00000000";
		ram_buffer(13272) := X"00000000";
		ram_buffer(13273) := X"00000000";
		ram_buffer(13274) := X"00000000";
		ram_buffer(13275) := X"00000000";
		ram_buffer(13276) := X"00000000";
		ram_buffer(13277) := X"00000000";
		ram_buffer(13278) := X"00000000";
		ram_buffer(13279) := X"00000000";
		ram_buffer(13280) := X"00000000";
		ram_buffer(13281) := X"00000000";
		ram_buffer(13282) := X"00000000";
		ram_buffer(13283) := X"00000000";
		ram_buffer(13284) := X"00000000";
		ram_buffer(13285) := X"00000000";
		ram_buffer(13286) := X"00000000";
		ram_buffer(13287) := X"00000000";
		ram_buffer(13288) := X"00000000";
		ram_buffer(13289) := X"00000000";
		ram_buffer(13290) := X"00000000";
		ram_buffer(13291) := X"00000000";
		ram_buffer(13292) := X"00000000";
		ram_buffer(13293) := X"00000000";
		ram_buffer(13294) := X"00000000";
		ram_buffer(13295) := X"00000000";
		ram_buffer(13296) := X"00000000";
		ram_buffer(13297) := X"00000000";
		ram_buffer(13298) := X"00000000";
		ram_buffer(13299) := X"00000000";
		ram_buffer(13300) := X"00000000";
		ram_buffer(13301) := X"00000000";
		ram_buffer(13302) := X"00000000";
		ram_buffer(13303) := X"00000000";
		ram_buffer(13304) := X"00000000";
		ram_buffer(13305) := X"00000000";
		ram_buffer(13306) := X"00000000";
		ram_buffer(13307) := X"00000000";
		ram_buffer(13308) := X"00000000";
		ram_buffer(13309) := X"00000000";
		ram_buffer(13310) := X"00000000";
		ram_buffer(13311) := X"00000000";
		ram_buffer(13312) := X"00000000";
		ram_buffer(13313) := X"00000000";
		ram_buffer(13314) := X"00000000";
		ram_buffer(13315) := X"00000000";
		ram_buffer(13316) := X"00000000";
		ram_buffer(13317) := X"00000000";
		ram_buffer(13318) := X"00000000";
		ram_buffer(13319) := X"00000000";
		ram_buffer(13320) := X"00000000";
		ram_buffer(13321) := X"00000000";
		ram_buffer(13322) := X"00000000";
		ram_buffer(13323) := X"00000000";
		ram_buffer(13324) := X"00000000";
		ram_buffer(13325) := X"00000000";
		ram_buffer(13326) := X"00000000";
		ram_buffer(13327) := X"00000000";
		ram_buffer(13328) := X"00000000";
		ram_buffer(13329) := X"00000000";
		ram_buffer(13330) := X"00000000";
		ram_buffer(13331) := X"00000000";
		ram_buffer(13332) := X"00000000";
		ram_buffer(13333) := X"00000000";
		ram_buffer(13334) := X"00000000";
		ram_buffer(13335) := X"00000000";
		ram_buffer(13336) := X"00000000";
		ram_buffer(13337) := X"00000000";
		ram_buffer(13338) := X"00000000";
		ram_buffer(13339) := X"00000000";
		ram_buffer(13340) := X"00000000";
		ram_buffer(13341) := X"00000000";
		ram_buffer(13342) := X"00000000";
		ram_buffer(13343) := X"00000000";
		ram_buffer(13344) := X"00000000";
		ram_buffer(13345) := X"00000000";
		ram_buffer(13346) := X"00000000";
		ram_buffer(13347) := X"00000000";
		ram_buffer(13348) := X"00000000";
		ram_buffer(13349) := X"00000000";
		ram_buffer(13350) := X"00000000";
		ram_buffer(13351) := X"00000000";
		ram_buffer(13352) := X"00000000";
		ram_buffer(13353) := X"00000000";
		ram_buffer(13354) := X"00000000";
		ram_buffer(13355) := X"00000000";
		ram_buffer(13356) := X"00000000";
		ram_buffer(13357) := X"00000000";
		ram_buffer(13358) := X"00000000";
		ram_buffer(13359) := X"00000000";
		ram_buffer(13360) := X"00000000";
		ram_buffer(13361) := X"00000000";
		ram_buffer(13362) := X"00000000";
		ram_buffer(13363) := X"00000000";
		ram_buffer(13364) := X"00000000";
		ram_buffer(13365) := X"00000000";
		ram_buffer(13366) := X"00000000";
		ram_buffer(13367) := X"00000000";
		ram_buffer(13368) := X"00000000";
		ram_buffer(13369) := X"00000000";
		ram_buffer(13370) := X"00000000";
		ram_buffer(13371) := X"00000000";
		ram_buffer(13372) := X"00000000";
		ram_buffer(13373) := X"00000000";
		ram_buffer(13374) := X"00000000";
		ram_buffer(13375) := X"00000000";
		ram_buffer(13376) := X"00000000";
		ram_buffer(13377) := X"00000000";
		ram_buffer(13378) := X"00000000";
		ram_buffer(13379) := X"00000000";
		ram_buffer(13380) := X"00000000";
		ram_buffer(13381) := X"00000000";
		ram_buffer(13382) := X"00000000";
		ram_buffer(13383) := X"00000000";
		ram_buffer(13384) := X"00000000";
		ram_buffer(13385) := X"00000000";
		ram_buffer(13386) := X"00000000";
		ram_buffer(13387) := X"00000000";
		ram_buffer(13388) := X"00000000";
		ram_buffer(13389) := X"00000000";
		ram_buffer(13390) := X"00000000";
		ram_buffer(13391) := X"00000000";
		ram_buffer(13392) := X"00000000";
		ram_buffer(13393) := X"00000000";
		ram_buffer(13394) := X"00000000";
		ram_buffer(13395) := X"00000000";
		ram_buffer(13396) := X"00000000";
		ram_buffer(13397) := X"00000000";
		ram_buffer(13398) := X"00000000";
		ram_buffer(13399) := X"00000000";
		ram_buffer(13400) := X"00000000";
		ram_buffer(13401) := X"00000000";
		ram_buffer(13402) := X"00000000";
		ram_buffer(13403) := X"00000000";
		ram_buffer(13404) := X"00000000";
		ram_buffer(13405) := X"00000000";
		ram_buffer(13406) := X"00000000";
		ram_buffer(13407) := X"00000000";
		ram_buffer(13408) := X"00000000";
		ram_buffer(13409) := X"00000000";
		ram_buffer(13410) := X"00000000";
		ram_buffer(13411) := X"00000000";
		ram_buffer(13412) := X"00000000";
		ram_buffer(13413) := X"00000000";
		ram_buffer(13414) := X"00000000";
		ram_buffer(13415) := X"00000000";
		ram_buffer(13416) := X"00000000";
		ram_buffer(13417) := X"00000000";
		ram_buffer(13418) := X"00000000";
		ram_buffer(13419) := X"00000000";
		ram_buffer(13420) := X"00000000";
		ram_buffer(13421) := X"00000000";
		ram_buffer(13422) := X"00000000";
		ram_buffer(13423) := X"00000000";
		ram_buffer(13424) := X"00000000";
		ram_buffer(13425) := X"00000000";
		ram_buffer(13426) := X"00000000";
		ram_buffer(13427) := X"00000000";
		ram_buffer(13428) := X"00000000";
		ram_buffer(13429) := X"00000000";
		ram_buffer(13430) := X"00000000";
		ram_buffer(13431) := X"00000000";
		ram_buffer(13432) := X"00000000";
		ram_buffer(13433) := X"00000000";
		ram_buffer(13434) := X"00000000";
		ram_buffer(13435) := X"00000000";
		ram_buffer(13436) := X"00000000";
		ram_buffer(13437) := X"00000000";
		ram_buffer(13438) := X"00000000";
		ram_buffer(13439) := X"00000000";
		ram_buffer(13440) := X"00000000";
		ram_buffer(13441) := X"00000000";
		ram_buffer(13442) := X"00000000";
		ram_buffer(13443) := X"00000000";
		ram_buffer(13444) := X"00000000";
		ram_buffer(13445) := X"00000000";
		ram_buffer(13446) := X"00000000";
		ram_buffer(13447) := X"00000000";
		ram_buffer(13448) := X"00000000";
		ram_buffer(13449) := X"00000000";
		ram_buffer(13450) := X"00000000";
		ram_buffer(13451) := X"00000000";
		ram_buffer(13452) := X"00000000";
		ram_buffer(13453) := X"00000000";
		ram_buffer(13454) := X"00000000";
		ram_buffer(13455) := X"00000000";
		ram_buffer(13456) := X"00000000";
		ram_buffer(13457) := X"00000000";
		ram_buffer(13458) := X"00000000";
		ram_buffer(13459) := X"00000000";
		ram_buffer(13460) := X"00000000";
		ram_buffer(13461) := X"00000000";
		ram_buffer(13462) := X"00000000";
		ram_buffer(13463) := X"00000000";
		ram_buffer(13464) := X"00000000";
		ram_buffer(13465) := X"00000000";
		ram_buffer(13466) := X"00000000";
		ram_buffer(13467) := X"00000000";
		ram_buffer(13468) := X"00000000";
		ram_buffer(13469) := X"00000000";
		ram_buffer(13470) := X"00000000";
		ram_buffer(13471) := X"00000000";
		ram_buffer(13472) := X"00000000";
		ram_buffer(13473) := X"00000000";
		ram_buffer(13474) := X"00000000";
		ram_buffer(13475) := X"00000000";
		ram_buffer(13476) := X"00000000";
		ram_buffer(13477) := X"00000000";
		ram_buffer(13478) := X"00000000";
		ram_buffer(13479) := X"00000000";
		ram_buffer(13480) := X"00000000";
		ram_buffer(13481) := X"00000000";
		ram_buffer(13482) := X"00000000";
		ram_buffer(13483) := X"00000000";
		ram_buffer(13484) := X"00000000";
		ram_buffer(13485) := X"00000000";
		ram_buffer(13486) := X"00000000";
		ram_buffer(13487) := X"00000000";
		ram_buffer(13488) := X"00000000";
		ram_buffer(13489) := X"00000000";
		ram_buffer(13490) := X"00000000";
		ram_buffer(13491) := X"00000000";
		ram_buffer(13492) := X"00000000";
		ram_buffer(13493) := X"00000000";
		ram_buffer(13494) := X"00000000";
		ram_buffer(13495) := X"00000000";
		ram_buffer(13496) := X"00000000";
		ram_buffer(13497) := X"00000000";
		ram_buffer(13498) := X"00000000";
		ram_buffer(13499) := X"00000000";
		ram_buffer(13500) := X"00000000";
		ram_buffer(13501) := X"00000000";
		ram_buffer(13502) := X"00000000";
		ram_buffer(13503) := X"00000000";
		ram_buffer(13504) := X"00000000";
		ram_buffer(13505) := X"00000000";
		ram_buffer(13506) := X"00000000";
		ram_buffer(13507) := X"00000000";
		ram_buffer(13508) := X"00000000";
		ram_buffer(13509) := X"00000000";
		ram_buffer(13510) := X"00000000";
		ram_buffer(13511) := X"00000000";
		ram_buffer(13512) := X"00000000";
		ram_buffer(13513) := X"00000000";
		ram_buffer(13514) := X"00000000";
		ram_buffer(13515) := X"00000000";
		ram_buffer(13516) := X"00000000";
		ram_buffer(13517) := X"00000000";
		ram_buffer(13518) := X"00000000";
		ram_buffer(13519) := X"00000000";
		ram_buffer(13520) := X"00000000";
		ram_buffer(13521) := X"00000000";
		ram_buffer(13522) := X"00000000";
		ram_buffer(13523) := X"00000000";
		ram_buffer(13524) := X"00000000";
		ram_buffer(13525) := X"00000000";
		ram_buffer(13526) := X"00000000";
		ram_buffer(13527) := X"00000000";
		ram_buffer(13528) := X"00000000";
		ram_buffer(13529) := X"00000000";
		ram_buffer(13530) := X"00000000";
		ram_buffer(13531) := X"00000000";
		ram_buffer(13532) := X"00000000";
		ram_buffer(13533) := X"00000000";
		ram_buffer(13534) := X"00000000";
		ram_buffer(13535) := X"00000000";
		ram_buffer(13536) := X"00000000";
		ram_buffer(13537) := X"00000000";
		ram_buffer(13538) := X"00000000";
		ram_buffer(13539) := X"00000000";
		ram_buffer(13540) := X"00000000";
		ram_buffer(13541) := X"00000000";
		ram_buffer(13542) := X"00000000";
		ram_buffer(13543) := X"00000000";
		ram_buffer(13544) := X"00000000";
		ram_buffer(13545) := X"00000000";
		ram_buffer(13546) := X"00000000";
		ram_buffer(13547) := X"00000000";
		ram_buffer(13548) := X"00000000";
		ram_buffer(13549) := X"00000000";
		ram_buffer(13550) := X"00000000";
		ram_buffer(13551) := X"00000000";
		ram_buffer(13552) := X"00000000";
		ram_buffer(13553) := X"00000000";
		ram_buffer(13554) := X"00000000";
		ram_buffer(13555) := X"00000000";
		ram_buffer(13556) := X"00000000";
		ram_buffer(13557) := X"00000000";
		ram_buffer(13558) := X"00000000";
		ram_buffer(13559) := X"00000000";
		ram_buffer(13560) := X"00000000";
		ram_buffer(13561) := X"00000000";
		ram_buffer(13562) := X"00000000";
		ram_buffer(13563) := X"00000000";
		ram_buffer(13564) := X"00000000";
		ram_buffer(13565) := X"00000000";
		ram_buffer(13566) := X"00000000";
		ram_buffer(13567) := X"00000000";
		ram_buffer(13568) := X"00000000";
		ram_buffer(13569) := X"00000000";
		ram_buffer(13570) := X"00000000";
		ram_buffer(13571) := X"00000000";
		ram_buffer(13572) := X"00000000";
		ram_buffer(13573) := X"00000000";
		ram_buffer(13574) := X"00000000";
		ram_buffer(13575) := X"00000000";
		ram_buffer(13576) := X"00000000";
		ram_buffer(13577) := X"00000000";
		ram_buffer(13578) := X"00000000";
		ram_buffer(13579) := X"00000000";
		ram_buffer(13580) := X"00000000";
		ram_buffer(13581) := X"00000000";
		ram_buffer(13582) := X"00000000";
		ram_buffer(13583) := X"00000000";
		ram_buffer(13584) := X"00000000";
		ram_buffer(13585) := X"00000000";
		ram_buffer(13586) := X"00000000";
		ram_buffer(13587) := X"00000000";
		ram_buffer(13588) := X"00000000";
		ram_buffer(13589) := X"00000000";
		ram_buffer(13590) := X"00000000";
		ram_buffer(13591) := X"00000000";
		ram_buffer(13592) := X"00000000";
		ram_buffer(13593) := X"00000000";
		ram_buffer(13594) := X"00000000";
		ram_buffer(13595) := X"00000000";
		ram_buffer(13596) := X"00000000";
		ram_buffer(13597) := X"00000000";
		ram_buffer(13598) := X"00000000";
		ram_buffer(13599) := X"00000000";
		ram_buffer(13600) := X"00000000";
		ram_buffer(13601) := X"00000000";
		ram_buffer(13602) := X"00000000";
		ram_buffer(13603) := X"00000000";
		ram_buffer(13604) := X"00000000";
		ram_buffer(13605) := X"00000000";
		ram_buffer(13606) := X"00000000";
		ram_buffer(13607) := X"00000000";
		ram_buffer(13608) := X"00000000";
		ram_buffer(13609) := X"00000000";
		ram_buffer(13610) := X"00000000";
		ram_buffer(13611) := X"00000000";
		ram_buffer(13612) := X"00000000";
		ram_buffer(13613) := X"00000000";
		ram_buffer(13614) := X"00000000";
		ram_buffer(13615) := X"00000000";
		ram_buffer(13616) := X"00000000";
		ram_buffer(13617) := X"00000000";
		ram_buffer(13618) := X"00000000";
		ram_buffer(13619) := X"00000000";
		ram_buffer(13620) := X"00000000";
		ram_buffer(13621) := X"00000000";
		ram_buffer(13622) := X"00000000";
		ram_buffer(13623) := X"00000000";
		ram_buffer(13624) := X"00000000";
		ram_buffer(13625) := X"00000000";
		ram_buffer(13626) := X"00000000";
		ram_buffer(13627) := X"00000000";
		ram_buffer(13628) := X"00000000";
		ram_buffer(13629) := X"00000000";
		ram_buffer(13630) := X"00000000";
		ram_buffer(13631) := X"00000000";
		ram_buffer(13632) := X"00000000";
		ram_buffer(13633) := X"00000000";
		ram_buffer(13634) := X"00000000";
		ram_buffer(13635) := X"00000000";
		ram_buffer(13636) := X"00000000";
		ram_buffer(13637) := X"00000000";
		ram_buffer(13638) := X"00000000";
		ram_buffer(13639) := X"00000000";
		ram_buffer(13640) := X"00000000";
		ram_buffer(13641) := X"00000000";
		ram_buffer(13642) := X"00000000";
		ram_buffer(13643) := X"00000000";
		ram_buffer(13644) := X"00000000";
		ram_buffer(13645) := X"00000000";
		ram_buffer(13646) := X"00000000";
		ram_buffer(13647) := X"00000000";
		ram_buffer(13648) := X"00000000";
		ram_buffer(13649) := X"00000000";
		ram_buffer(13650) := X"00000000";
		ram_buffer(13651) := X"00000000";
		ram_buffer(13652) := X"00000000";
		ram_buffer(13653) := X"00000000";
		ram_buffer(13654) := X"00000000";
		ram_buffer(13655) := X"00000000";
		ram_buffer(13656) := X"00000000";
		ram_buffer(13657) := X"00000000";
		ram_buffer(13658) := X"00000000";
		ram_buffer(13659) := X"00000000";
		ram_buffer(13660) := X"00000000";
		ram_buffer(13661) := X"00000000";
		ram_buffer(13662) := X"00000000";
		ram_buffer(13663) := X"00000000";
		ram_buffer(13664) := X"00000000";
		ram_buffer(13665) := X"00000000";
		ram_buffer(13666) := X"00000000";
		ram_buffer(13667) := X"00000000";
		ram_buffer(13668) := X"00000000";
		ram_buffer(13669) := X"00000000";
		ram_buffer(13670) := X"00000000";
		ram_buffer(13671) := X"00000000";
		ram_buffer(13672) := X"00000000";
		ram_buffer(13673) := X"00000000";
		ram_buffer(13674) := X"00000000";
		ram_buffer(13675) := X"00000000";
		ram_buffer(13676) := X"00000000";
		ram_buffer(13677) := X"00000000";
		ram_buffer(13678) := X"00000000";
		ram_buffer(13679) := X"00000000";
		ram_buffer(13680) := X"00000000";
		ram_buffer(13681) := X"00000000";
		ram_buffer(13682) := X"00000000";
		ram_buffer(13683) := X"00000000";
		ram_buffer(13684) := X"00000000";
		ram_buffer(13685) := X"00000000";
		ram_buffer(13686) := X"00000000";
		ram_buffer(13687) := X"00000000";
		ram_buffer(13688) := X"00000000";
		ram_buffer(13689) := X"00000000";
		ram_buffer(13690) := X"00000000";
		ram_buffer(13691) := X"00000000";
		ram_buffer(13692) := X"00000000";
		ram_buffer(13693) := X"00000000";
		ram_buffer(13694) := X"00000000";
		ram_buffer(13695) := X"00000000";
		ram_buffer(13696) := X"00000000";
		ram_buffer(13697) := X"00000000";
		ram_buffer(13698) := X"00000000";
		ram_buffer(13699) := X"00000000";
		ram_buffer(13700) := X"00000000";
		ram_buffer(13701) := X"00000000";
		ram_buffer(13702) := X"00000000";
		ram_buffer(13703) := X"00000000";
		ram_buffer(13704) := X"00000000";
		ram_buffer(13705) := X"00000000";
		ram_buffer(13706) := X"00000000";
		ram_buffer(13707) := X"00000000";
		ram_buffer(13708) := X"00000000";
		ram_buffer(13709) := X"00000000";
		ram_buffer(13710) := X"00000000";
		ram_buffer(13711) := X"00000000";
		ram_buffer(13712) := X"00000000";
		ram_buffer(13713) := X"00000000";
		ram_buffer(13714) := X"00000000";
		ram_buffer(13715) := X"00000000";
		ram_buffer(13716) := X"00000000";
		ram_buffer(13717) := X"00000000";
		ram_buffer(13718) := X"00000000";
		ram_buffer(13719) := X"00000000";
		ram_buffer(13720) := X"00000000";
		ram_buffer(13721) := X"00000000";
		ram_buffer(13722) := X"00000000";
		ram_buffer(13723) := X"00000000";
		ram_buffer(13724) := X"00000000";
		ram_buffer(13725) := X"00000000";
		ram_buffer(13726) := X"00000000";
		ram_buffer(13727) := X"00000000";
		ram_buffer(13728) := X"00000000";
		ram_buffer(13729) := X"00000000";
		ram_buffer(13730) := X"00000000";
		ram_buffer(13731) := X"00000000";
		ram_buffer(13732) := X"00000000";
		ram_buffer(13733) := X"00000000";
		ram_buffer(13734) := X"00000000";
		ram_buffer(13735) := X"00000000";
		ram_buffer(13736) := X"00000000";
		ram_buffer(13737) := X"00000000";
		ram_buffer(13738) := X"00000000";
		ram_buffer(13739) := X"00000000";
		ram_buffer(13740) := X"00000000";
		ram_buffer(13741) := X"00000000";
		ram_buffer(13742) := X"00000000";
		ram_buffer(13743) := X"00000000";
		ram_buffer(13744) := X"00000000";
		ram_buffer(13745) := X"00000000";
		ram_buffer(13746) := X"00000000";
		ram_buffer(13747) := X"00000000";
		ram_buffer(13748) := X"00000000";
		ram_buffer(13749) := X"00000000";
		ram_buffer(13750) := X"00000000";
		ram_buffer(13751) := X"00000000";
		ram_buffer(13752) := X"00000000";
		ram_buffer(13753) := X"00000000";
		ram_buffer(13754) := X"00000000";
		ram_buffer(13755) := X"00000000";
		ram_buffer(13756) := X"00000000";
		ram_buffer(13757) := X"00000000";
		ram_buffer(13758) := X"00000000";
		ram_buffer(13759) := X"00000000";
		ram_buffer(13760) := X"00000000";
		ram_buffer(13761) := X"00000000";
		ram_buffer(13762) := X"00000000";
		ram_buffer(13763) := X"00000000";
		ram_buffer(13764) := X"00000000";
		ram_buffer(13765) := X"00000000";
		ram_buffer(13766) := X"00000000";
		ram_buffer(13767) := X"00000000";
		ram_buffer(13768) := X"00000000";
		ram_buffer(13769) := X"00000000";
		ram_buffer(13770) := X"00000000";
		ram_buffer(13771) := X"00000000";
		ram_buffer(13772) := X"00000000";
		ram_buffer(13773) := X"00000000";
		ram_buffer(13774) := X"00000000";
		ram_buffer(13775) := X"00000000";
		ram_buffer(13776) := X"00000000";
		ram_buffer(13777) := X"00000000";
		ram_buffer(13778) := X"00000000";
		ram_buffer(13779) := X"00000000";
		ram_buffer(13780) := X"00000000";
		ram_buffer(13781) := X"00000000";
		ram_buffer(13782) := X"00000000";
		ram_buffer(13783) := X"00000000";
		ram_buffer(13784) := X"00000000";
		ram_buffer(13785) := X"00000000";
		ram_buffer(13786) := X"00000000";
		ram_buffer(13787) := X"00000000";
		ram_buffer(13788) := X"00000000";
		ram_buffer(13789) := X"00000000";
		ram_buffer(13790) := X"00000000";
		ram_buffer(13791) := X"00000000";
		ram_buffer(13792) := X"00000000";
		ram_buffer(13793) := X"00000000";
		ram_buffer(13794) := X"00000000";
		ram_buffer(13795) := X"00000000";
		ram_buffer(13796) := X"00000000";
		ram_buffer(13797) := X"00000000";
		ram_buffer(13798) := X"00000000";
		ram_buffer(13799) := X"00000000";
		ram_buffer(13800) := X"00000000";
		ram_buffer(13801) := X"00000000";
		ram_buffer(13802) := X"00000000";
		ram_buffer(13803) := X"00000000";
		ram_buffer(13804) := X"00000000";
		ram_buffer(13805) := X"00000000";
		ram_buffer(13806) := X"00000000";
		ram_buffer(13807) := X"00000000";
		ram_buffer(13808) := X"00000000";
		ram_buffer(13809) := X"00000000";
		ram_buffer(13810) := X"00000000";
		ram_buffer(13811) := X"00000000";
		ram_buffer(13812) := X"00000000";
		ram_buffer(13813) := X"00000000";
		ram_buffer(13814) := X"00000000";
		ram_buffer(13815) := X"00000000";
		ram_buffer(13816) := X"00000000";
		ram_buffer(13817) := X"00000000";
		ram_buffer(13818) := X"00000000";
		ram_buffer(13819) := X"00000000";
		ram_buffer(13820) := X"00000000";
		ram_buffer(13821) := X"00000000";
		ram_buffer(13822) := X"00000000";
		ram_buffer(13823) := X"00000000";
		ram_buffer(13824) := X"00000000";
		ram_buffer(13825) := X"00000000";
		ram_buffer(13826) := X"00000000";
		ram_buffer(13827) := X"00000000";
		ram_buffer(13828) := X"00000000";
		ram_buffer(13829) := X"00000000";
		ram_buffer(13830) := X"00000000";
		ram_buffer(13831) := X"00000000";
		ram_buffer(13832) := X"00000000";
		ram_buffer(13833) := X"00000000";
		ram_buffer(13834) := X"00000000";
		ram_buffer(13835) := X"00000000";
		ram_buffer(13836) := X"00000000";
		ram_buffer(13837) := X"00000000";
		ram_buffer(13838) := X"00000000";
		ram_buffer(13839) := X"00000000";
		ram_buffer(13840) := X"00000000";
		ram_buffer(13841) := X"00000000";
		ram_buffer(13842) := X"00000000";
		ram_buffer(13843) := X"00000000";
		ram_buffer(13844) := X"00000000";
		ram_buffer(13845) := X"00000000";
		ram_buffer(13846) := X"00000000";
		ram_buffer(13847) := X"00000000";
		ram_buffer(13848) := X"00000000";
		ram_buffer(13849) := X"00000000";
		ram_buffer(13850) := X"00000000";
		ram_buffer(13851) := X"00000000";
		ram_buffer(13852) := X"00000000";
		ram_buffer(13853) := X"00000000";
		ram_buffer(13854) := X"00000000";
		ram_buffer(13855) := X"00000000";
		ram_buffer(13856) := X"00000000";
		ram_buffer(13857) := X"00000000";
		ram_buffer(13858) := X"00000000";
		ram_buffer(13859) := X"00000000";
		ram_buffer(13860) := X"00000000";
		ram_buffer(13861) := X"00000000";
		ram_buffer(13862) := X"00000000";
		ram_buffer(13863) := X"00000000";
		ram_buffer(13864) := X"00000000";
		ram_buffer(13865) := X"00000000";
		ram_buffer(13866) := X"00000000";
		ram_buffer(13867) := X"00000000";
		ram_buffer(13868) := X"00000000";
		ram_buffer(13869) := X"00000000";
		ram_buffer(13870) := X"00000000";
		ram_buffer(13871) := X"00000000";
		ram_buffer(13872) := X"00000000";
		ram_buffer(13873) := X"00000000";
		ram_buffer(13874) := X"00000000";
		ram_buffer(13875) := X"00000000";
		ram_buffer(13876) := X"00000000";
		ram_buffer(13877) := X"00000000";
		ram_buffer(13878) := X"00000000";
		ram_buffer(13879) := X"00000000";
		ram_buffer(13880) := X"00000000";
		ram_buffer(13881) := X"00000000";
		ram_buffer(13882) := X"00000000";
		ram_buffer(13883) := X"00000000";
		ram_buffer(13884) := X"00000000";
		ram_buffer(13885) := X"00000000";
		ram_buffer(13886) := X"00000000";
		ram_buffer(13887) := X"00000000";
		ram_buffer(13888) := X"00000000";
		ram_buffer(13889) := X"00000000";
		ram_buffer(13890) := X"00000000";
		ram_buffer(13891) := X"00000000";
		ram_buffer(13892) := X"00000000";
		ram_buffer(13893) := X"00000000";
		ram_buffer(13894) := X"00000000";
		ram_buffer(13895) := X"00000000";
		ram_buffer(13896) := X"00000000";
		ram_buffer(13897) := X"00000000";
		ram_buffer(13898) := X"00000000";
		ram_buffer(13899) := X"00000000";
		ram_buffer(13900) := X"00000000";
		ram_buffer(13901) := X"00000000";
		ram_buffer(13902) := X"00000000";
		ram_buffer(13903) := X"00000000";
		ram_buffer(13904) := X"00000000";
		ram_buffer(13905) := X"00000000";
		ram_buffer(13906) := X"00000000";
		ram_buffer(13907) := X"00000000";
		ram_buffer(13908) := X"00000000";
		ram_buffer(13909) := X"00000000";
		ram_buffer(13910) := X"00000000";
		ram_buffer(13911) := X"00000000";
		ram_buffer(13912) := X"00000000";
		ram_buffer(13913) := X"00000000";
		ram_buffer(13914) := X"00000000";
		ram_buffer(13915) := X"00000000";
		ram_buffer(13916) := X"00000000";
		ram_buffer(13917) := X"00000000";
		ram_buffer(13918) := X"00000000";
		ram_buffer(13919) := X"00000000";
		ram_buffer(13920) := X"00000000";
		ram_buffer(13921) := X"00000000";
		ram_buffer(13922) := X"00000000";
		ram_buffer(13923) := X"00000000";
		ram_buffer(13924) := X"00000000";
		ram_buffer(13925) := X"00000000";
		ram_buffer(13926) := X"00000000";
		ram_buffer(13927) := X"00000000";
		ram_buffer(13928) := X"00000000";
		ram_buffer(13929) := X"00000000";
		ram_buffer(13930) := X"00000000";
		ram_buffer(13931) := X"00000000";
		ram_buffer(13932) := X"00000000";
		ram_buffer(13933) := X"00000000";
		ram_buffer(13934) := X"00000000";
		ram_buffer(13935) := X"00000000";
		ram_buffer(13936) := X"00000000";
		ram_buffer(13937) := X"00000000";
		ram_buffer(13938) := X"00000000";
		ram_buffer(13939) := X"00000000";
		ram_buffer(13940) := X"00000000";
		ram_buffer(13941) := X"00000000";
		ram_buffer(13942) := X"00000000";
		ram_buffer(13943) := X"00000000";
		ram_buffer(13944) := X"00000000";
		ram_buffer(13945) := X"00000000";
		ram_buffer(13946) := X"00000000";
		ram_buffer(13947) := X"00000000";
		ram_buffer(13948) := X"00000000";
		ram_buffer(13949) := X"00000000";
		ram_buffer(13950) := X"00000000";
		ram_buffer(13951) := X"00000000";
		ram_buffer(13952) := X"00000000";
		ram_buffer(13953) := X"00000000";
		ram_buffer(13954) := X"00000000";
		ram_buffer(13955) := X"00000000";
		ram_buffer(13956) := X"00000000";
		ram_buffer(13957) := X"00000000";
		ram_buffer(13958) := X"00000000";
		ram_buffer(13959) := X"00000000";
		ram_buffer(13960) := X"00000000";
		ram_buffer(13961) := X"00000000";
		ram_buffer(13962) := X"00000000";
		ram_buffer(13963) := X"00000000";
		ram_buffer(13964) := X"00000000";
		ram_buffer(13965) := X"00000000";
		ram_buffer(13966) := X"00000000";
		ram_buffer(13967) := X"00000000";
		ram_buffer(13968) := X"00000000";
		ram_buffer(13969) := X"00000000";
		ram_buffer(13970) := X"00000000";
		ram_buffer(13971) := X"00000000";
		ram_buffer(13972) := X"00000000";
		ram_buffer(13973) := X"00000000";
		ram_buffer(13974) := X"00000000";
		ram_buffer(13975) := X"00000000";
		ram_buffer(13976) := X"00000000";
		ram_buffer(13977) := X"00000000";
		ram_buffer(13978) := X"00000000";
		ram_buffer(13979) := X"00000000";
		ram_buffer(13980) := X"00000000";
		ram_buffer(13981) := X"00000000";
		ram_buffer(13982) := X"00000000";
		ram_buffer(13983) := X"00000000";
		ram_buffer(13984) := X"00000000";
		ram_buffer(13985) := X"00000000";
		ram_buffer(13986) := X"00000000";
		ram_buffer(13987) := X"00000000";
		ram_buffer(13988) := X"00000000";
		ram_buffer(13989) := X"00000000";
		ram_buffer(13990) := X"00000000";
		ram_buffer(13991) := X"00000000";
		ram_buffer(13992) := X"00000000";
		ram_buffer(13993) := X"00000000";
		ram_buffer(13994) := X"00000000";
		ram_buffer(13995) := X"00000000";
		ram_buffer(13996) := X"00000000";
		ram_buffer(13997) := X"00000000";
		ram_buffer(13998) := X"00000000";
		ram_buffer(13999) := X"00000000";
		ram_buffer(14000) := X"00000000";
		ram_buffer(14001) := X"00000000";
		ram_buffer(14002) := X"00000000";
		ram_buffer(14003) := X"00000000";
		ram_buffer(14004) := X"00000000";
		ram_buffer(14005) := X"00000000";
		ram_buffer(14006) := X"00000000";
		ram_buffer(14007) := X"00000000";
		ram_buffer(14008) := X"00000000";
		ram_buffer(14009) := X"00000000";
		ram_buffer(14010) := X"00000000";
		ram_buffer(14011) := X"00000000";
		ram_buffer(14012) := X"00000000";
		ram_buffer(14013) := X"00000000";
		ram_buffer(14014) := X"00000000";
		ram_buffer(14015) := X"00000000";
		ram_buffer(14016) := X"00000000";
		ram_buffer(14017) := X"00000000";
		ram_buffer(14018) := X"00000000";
		ram_buffer(14019) := X"00000000";
		ram_buffer(14020) := X"00000000";
		ram_buffer(14021) := X"00000000";
		ram_buffer(14022) := X"00000000";
		ram_buffer(14023) := X"00000000";
		ram_buffer(14024) := X"00000000";
		ram_buffer(14025) := X"00000000";
		ram_buffer(14026) := X"00000000";
		ram_buffer(14027) := X"00000000";
		ram_buffer(14028) := X"00000000";
		ram_buffer(14029) := X"00000000";
		ram_buffer(14030) := X"00000000";
		ram_buffer(14031) := X"00000000";
		ram_buffer(14032) := X"00000000";
		ram_buffer(14033) := X"00000000";
		ram_buffer(14034) := X"00000000";
		ram_buffer(14035) := X"00000000";
		ram_buffer(14036) := X"00000000";
		ram_buffer(14037) := X"00000000";
		ram_buffer(14038) := X"00000000";
		ram_buffer(14039) := X"00000000";
		ram_buffer(14040) := X"00000000";
		ram_buffer(14041) := X"00000000";
		ram_buffer(14042) := X"00000000";
		ram_buffer(14043) := X"00000000";
		ram_buffer(14044) := X"00000000";
		ram_buffer(14045) := X"00000000";
		ram_buffer(14046) := X"00000000";
		ram_buffer(14047) := X"00000000";
		ram_buffer(14048) := X"00000000";
		ram_buffer(14049) := X"00000000";
		ram_buffer(14050) := X"00000000";
		ram_buffer(14051) := X"00000000";
		ram_buffer(14052) := X"00000000";
		ram_buffer(14053) := X"00000000";
		ram_buffer(14054) := X"00000000";
		ram_buffer(14055) := X"00000000";
		ram_buffer(14056) := X"00000000";
		ram_buffer(14057) := X"00000000";
		ram_buffer(14058) := X"00000000";
		ram_buffer(14059) := X"00000000";
		ram_buffer(14060) := X"00000000";
		ram_buffer(14061) := X"00000000";
		ram_buffer(14062) := X"00000000";
		ram_buffer(14063) := X"00000000";
		ram_buffer(14064) := X"00000000";
		ram_buffer(14065) := X"00000000";
		ram_buffer(14066) := X"00000000";
		ram_buffer(14067) := X"00000000";
		ram_buffer(14068) := X"00000000";
		ram_buffer(14069) := X"00000000";
		ram_buffer(14070) := X"00000000";
		ram_buffer(14071) := X"00000000";
		ram_buffer(14072) := X"00000000";
		ram_buffer(14073) := X"00000000";
		ram_buffer(14074) := X"00000000";
		ram_buffer(14075) := X"00000000";
		ram_buffer(14076) := X"00000000";
		ram_buffer(14077) := X"00000000";
		ram_buffer(14078) := X"00000000";
		ram_buffer(14079) := X"00000000";
		ram_buffer(14080) := X"00000000";
		ram_buffer(14081) := X"00000000";
		ram_buffer(14082) := X"00000000";
		ram_buffer(14083) := X"00000000";
		ram_buffer(14084) := X"00000000";
		ram_buffer(14085) := X"00000000";
		ram_buffer(14086) := X"00000000";
		ram_buffer(14087) := X"00000000";
		ram_buffer(14088) := X"00000000";
		ram_buffer(14089) := X"00000000";
		ram_buffer(14090) := X"00000000";
		ram_buffer(14091) := X"00000000";
		ram_buffer(14092) := X"00000000";
		ram_buffer(14093) := X"00000000";
		ram_buffer(14094) := X"00000000";
		ram_buffer(14095) := X"00000000";
		ram_buffer(14096) := X"00000000";
		ram_buffer(14097) := X"00000000";
		ram_buffer(14098) := X"00000000";
		ram_buffer(14099) := X"00000000";
		ram_buffer(14100) := X"00000000";
		ram_buffer(14101) := X"00000000";
		ram_buffer(14102) := X"00000000";
		ram_buffer(14103) := X"00000000";
		ram_buffer(14104) := X"00000000";
		ram_buffer(14105) := X"00000000";
		ram_buffer(14106) := X"00000000";
		ram_buffer(14107) := X"00000000";
		ram_buffer(14108) := X"00000000";
		ram_buffer(14109) := X"00000000";
		ram_buffer(14110) := X"00000000";
		ram_buffer(14111) := X"00000000";
		ram_buffer(14112) := X"00000000";
		ram_buffer(14113) := X"00000000";
		ram_buffer(14114) := X"00000000";
		ram_buffer(14115) := X"00000000";
		ram_buffer(14116) := X"00000000";
		ram_buffer(14117) := X"00000000";
		ram_buffer(14118) := X"00000000";
		ram_buffer(14119) := X"00000000";
		ram_buffer(14120) := X"00000000";
		ram_buffer(14121) := X"00000000";
		ram_buffer(14122) := X"00000000";
		ram_buffer(14123) := X"00000000";
		ram_buffer(14124) := X"00000000";
		ram_buffer(14125) := X"00000000";
		ram_buffer(14126) := X"00000000";
		ram_buffer(14127) := X"00000000";
		ram_buffer(14128) := X"00000000";
		ram_buffer(14129) := X"00000000";
		ram_buffer(14130) := X"00000000";
		ram_buffer(14131) := X"00000000";
		ram_buffer(14132) := X"00000000";
		ram_buffer(14133) := X"00000000";
		ram_buffer(14134) := X"00000000";
		ram_buffer(14135) := X"00000000";
		ram_buffer(14136) := X"00000000";
		ram_buffer(14137) := X"00000000";
		ram_buffer(14138) := X"00000000";
		ram_buffer(14139) := X"00000000";
		ram_buffer(14140) := X"00000000";
		ram_buffer(14141) := X"00000000";
		ram_buffer(14142) := X"00000000";
		ram_buffer(14143) := X"00000000";
		ram_buffer(14144) := X"00000000";
		ram_buffer(14145) := X"00000000";
		ram_buffer(14146) := X"00000000";
		ram_buffer(14147) := X"00000000";
		ram_buffer(14148) := X"00000000";
		ram_buffer(14149) := X"00000000";
		ram_buffer(14150) := X"00000000";
		ram_buffer(14151) := X"00000000";
		ram_buffer(14152) := X"00000000";
		ram_buffer(14153) := X"00000000";
		ram_buffer(14154) := X"00000000";
		ram_buffer(14155) := X"00000000";
		ram_buffer(14156) := X"00000000";
		ram_buffer(14157) := X"00000000";
		ram_buffer(14158) := X"00000000";
		ram_buffer(14159) := X"00000000";
		ram_buffer(14160) := X"00000000";
		ram_buffer(14161) := X"00000000";
		ram_buffer(14162) := X"00000000";
		ram_buffer(14163) := X"00000000";
		ram_buffer(14164) := X"00000000";
		ram_buffer(14165) := X"00000000";
		ram_buffer(14166) := X"00000000";
		ram_buffer(14167) := X"00000000";
		ram_buffer(14168) := X"00000000";
		ram_buffer(14169) := X"00000000";
		ram_buffer(14170) := X"00000000";
		ram_buffer(14171) := X"00000000";
		ram_buffer(14172) := X"00000000";
		ram_buffer(14173) := X"00000000";
		ram_buffer(14174) := X"00000000";
		ram_buffer(14175) := X"00000000";
		ram_buffer(14176) := X"00000000";
		ram_buffer(14177) := X"00000000";
		ram_buffer(14178) := X"00000000";
		ram_buffer(14179) := X"00000000";
		ram_buffer(14180) := X"00000000";
		ram_buffer(14181) := X"00000000";
		ram_buffer(14182) := X"00000000";
		ram_buffer(14183) := X"00000000";
		ram_buffer(14184) := X"00000000";
		ram_buffer(14185) := X"00000000";
		ram_buffer(14186) := X"00000000";
		ram_buffer(14187) := X"00000000";
		ram_buffer(14188) := X"00000000";
		ram_buffer(14189) := X"00000000";
		ram_buffer(14190) := X"00000000";
		ram_buffer(14191) := X"00000000";
		ram_buffer(14192) := X"00000000";
		ram_buffer(14193) := X"00000000";
		ram_buffer(14194) := X"00000000";
		ram_buffer(14195) := X"00000000";
		ram_buffer(14196) := X"00000000";
		ram_buffer(14197) := X"00000000";
		ram_buffer(14198) := X"00000000";
		ram_buffer(14199) := X"00000000";
		ram_buffer(14200) := X"00000000";
		ram_buffer(14201) := X"00000000";
		ram_buffer(14202) := X"00000000";
		ram_buffer(14203) := X"00000000";
		ram_buffer(14204) := X"00000000";
		ram_buffer(14205) := X"00000000";
		ram_buffer(14206) := X"00000000";
		ram_buffer(14207) := X"00000000";
		ram_buffer(14208) := X"00000000";
		ram_buffer(14209) := X"00000000";
		ram_buffer(14210) := X"00000000";
		ram_buffer(14211) := X"00000000";
		ram_buffer(14212) := X"00000000";
		ram_buffer(14213) := X"00000000";
		ram_buffer(14214) := X"00000000";
		ram_buffer(14215) := X"00000000";
		ram_buffer(14216) := X"00000000";
		ram_buffer(14217) := X"00000000";
		ram_buffer(14218) := X"00000000";
		ram_buffer(14219) := X"00000000";
		ram_buffer(14220) := X"00000000";
		ram_buffer(14221) := X"00000000";
		ram_buffer(14222) := X"00000000";
		ram_buffer(14223) := X"00000000";
		ram_buffer(14224) := X"00000000";
		ram_buffer(14225) := X"00000000";
		ram_buffer(14226) := X"00000000";
		ram_buffer(14227) := X"00000000";
		ram_buffer(14228) := X"00000000";
		ram_buffer(14229) := X"00000000";
		ram_buffer(14230) := X"00000000";
		ram_buffer(14231) := X"00000000";
		ram_buffer(14232) := X"00000000";
		ram_buffer(14233) := X"00000000";
		ram_buffer(14234) := X"00000000";
		ram_buffer(14235) := X"00000000";
		ram_buffer(14236) := X"00000000";
		ram_buffer(14237) := X"00000000";
		ram_buffer(14238) := X"00000000";
		ram_buffer(14239) := X"00000000";
		ram_buffer(14240) := X"00000000";
		ram_buffer(14241) := X"00000000";
		ram_buffer(14242) := X"00000000";
		ram_buffer(14243) := X"00000000";
		ram_buffer(14244) := X"00000000";
		ram_buffer(14245) := X"00000000";
		ram_buffer(14246) := X"00000000";
		ram_buffer(14247) := X"00000000";
		ram_buffer(14248) := X"00000000";
		ram_buffer(14249) := X"00000000";
		ram_buffer(14250) := X"00000000";
		ram_buffer(14251) := X"00000000";
		ram_buffer(14252) := X"00000000";
		ram_buffer(14253) := X"00000000";
		ram_buffer(14254) := X"00000000";
		ram_buffer(14255) := X"00000000";
		ram_buffer(14256) := X"00000000";
		ram_buffer(14257) := X"00000000";
		ram_buffer(14258) := X"00000000";
		ram_buffer(14259) := X"00000000";
		ram_buffer(14260) := X"00000000";
		ram_buffer(14261) := X"00000000";
		ram_buffer(14262) := X"00000000";
		ram_buffer(14263) := X"00000000";
		ram_buffer(14264) := X"00000000";
		ram_buffer(14265) := X"00000000";
		ram_buffer(14266) := X"00000000";
		ram_buffer(14267) := X"00000000";
		ram_buffer(14268) := X"00000000";
		ram_buffer(14269) := X"00000000";
		ram_buffer(14270) := X"00000000";
		ram_buffer(14271) := X"00000000";
		ram_buffer(14272) := X"00000000";
		ram_buffer(14273) := X"00000000";
		ram_buffer(14274) := X"00000000";
		ram_buffer(14275) := X"00000000";
		ram_buffer(14276) := X"00000000";
		ram_buffer(14277) := X"00000000";
		ram_buffer(14278) := X"00000000";
		ram_buffer(14279) := X"00000000";
		ram_buffer(14280) := X"00000000";
		ram_buffer(14281) := X"00000000";
		ram_buffer(14282) := X"00000000";
		ram_buffer(14283) := X"00000000";
		ram_buffer(14284) := X"00000000";
		ram_buffer(14285) := X"00000000";
		ram_buffer(14286) := X"00000000";
		ram_buffer(14287) := X"00000000";
		ram_buffer(14288) := X"00000000";
		ram_buffer(14289) := X"00000000";
		ram_buffer(14290) := X"00000000";
		ram_buffer(14291) := X"00000000";
		ram_buffer(14292) := X"00000000";
		ram_buffer(14293) := X"00000000";
		ram_buffer(14294) := X"00000000";
		ram_buffer(14295) := X"00000000";
		ram_buffer(14296) := X"00000000";
		ram_buffer(14297) := X"00000000";
		ram_buffer(14298) := X"00000000";
		ram_buffer(14299) := X"00000000";
		ram_buffer(14300) := X"00000000";
		ram_buffer(14301) := X"00000000";
		ram_buffer(14302) := X"00000000";
		ram_buffer(14303) := X"00000000";
		ram_buffer(14304) := X"00000000";
		ram_buffer(14305) := X"00000000";
		ram_buffer(14306) := X"00000000";
		ram_buffer(14307) := X"00000000";
		ram_buffer(14308) := X"00000000";
		ram_buffer(14309) := X"00000000";
		ram_buffer(14310) := X"00000000";
		ram_buffer(14311) := X"00000000";
		ram_buffer(14312) := X"00000000";
		ram_buffer(14313) := X"00000000";
		ram_buffer(14314) := X"00000000";
		ram_buffer(14315) := X"00000000";
		ram_buffer(14316) := X"00000000";
		ram_buffer(14317) := X"00000000";
		ram_buffer(14318) := X"00000000";
		ram_buffer(14319) := X"00000000";
		ram_buffer(14320) := X"00000000";
		ram_buffer(14321) := X"00000000";
		ram_buffer(14322) := X"00000000";
		ram_buffer(14323) := X"00000000";
		ram_buffer(14324) := X"00000000";
		ram_buffer(14325) := X"00000000";
		ram_buffer(14326) := X"00000000";
		ram_buffer(14327) := X"00000000";
		ram_buffer(14328) := X"00000000";
		ram_buffer(14329) := X"00000000";
		ram_buffer(14330) := X"00000000";
		ram_buffer(14331) := X"00000000";
		ram_buffer(14332) := X"00000000";
		ram_buffer(14333) := X"00000000";
		ram_buffer(14334) := X"00000000";
		ram_buffer(14335) := X"00000000";
		ram_buffer(14336) := X"00000000";
		ram_buffer(14337) := X"00000000";
		ram_buffer(14338) := X"00000000";
		ram_buffer(14339) := X"00000000";
		ram_buffer(14340) := X"00000000";
		ram_buffer(14341) := X"00000000";
		ram_buffer(14342) := X"00000000";
		ram_buffer(14343) := X"00000000";
		ram_buffer(14344) := X"00000000";
		ram_buffer(14345) := X"00000000";
		ram_buffer(14346) := X"00000000";
		ram_buffer(14347) := X"00000000";
		ram_buffer(14348) := X"00000000";
		ram_buffer(14349) := X"00000000";
		ram_buffer(14350) := X"00000000";
		ram_buffer(14351) := X"00000000";
		ram_buffer(14352) := X"00000000";
		ram_buffer(14353) := X"00000000";
		ram_buffer(14354) := X"00000000";
		ram_buffer(14355) := X"00000000";
		ram_buffer(14356) := X"00000000";
		ram_buffer(14357) := X"00000000";
		ram_buffer(14358) := X"00000000";
		ram_buffer(14359) := X"00000000";
		ram_buffer(14360) := X"00000000";
		ram_buffer(14361) := X"00000000";
		ram_buffer(14362) := X"00000000";
		ram_buffer(14363) := X"00000000";
		ram_buffer(14364) := X"00000000";
		ram_buffer(14365) := X"00000000";
		ram_buffer(14366) := X"00000000";
		ram_buffer(14367) := X"00000000";
		ram_buffer(14368) := X"00000000";
		ram_buffer(14369) := X"00000000";
		ram_buffer(14370) := X"00000000";
		ram_buffer(14371) := X"00000000";
		ram_buffer(14372) := X"00000000";
		ram_buffer(14373) := X"00000000";
		ram_buffer(14374) := X"00000000";
		ram_buffer(14375) := X"00000000";
		ram_buffer(14376) := X"00000000";
		ram_buffer(14377) := X"00000000";
		ram_buffer(14378) := X"00000000";
		ram_buffer(14379) := X"00000000";
		ram_buffer(14380) := X"00000000";
		ram_buffer(14381) := X"00000000";
		ram_buffer(14382) := X"00000000";
		ram_buffer(14383) := X"00000000";
		ram_buffer(14384) := X"00000000";
		ram_buffer(14385) := X"00000000";
		ram_buffer(14386) := X"00000000";
		ram_buffer(14387) := X"00000000";
		ram_buffer(14388) := X"00000000";
		ram_buffer(14389) := X"00000000";
		ram_buffer(14390) := X"00000000";
		ram_buffer(14391) := X"00000000";
		ram_buffer(14392) := X"00000000";
		ram_buffer(14393) := X"00000000";
		ram_buffer(14394) := X"00000000";
		ram_buffer(14395) := X"00000000";
		ram_buffer(14396) := X"00000000";
		ram_buffer(14397) := X"00000000";
		ram_buffer(14398) := X"00000000";
		ram_buffer(14399) := X"00000000";
		ram_buffer(14400) := X"00000000";
		ram_buffer(14401) := X"00000000";
		ram_buffer(14402) := X"00000000";
		ram_buffer(14403) := X"00000000";
		ram_buffer(14404) := X"00000000";
		ram_buffer(14405) := X"00000000";
		ram_buffer(14406) := X"00000000";
		ram_buffer(14407) := X"00000000";
		ram_buffer(14408) := X"00000000";
		ram_buffer(14409) := X"00000000";
		ram_buffer(14410) := X"00000000";
		ram_buffer(14411) := X"00000000";
		ram_buffer(14412) := X"00000000";
		ram_buffer(14413) := X"00000000";
		ram_buffer(14414) := X"00000000";
		ram_buffer(14415) := X"00000000";
		ram_buffer(14416) := X"00000000";
		ram_buffer(14417) := X"00000000";
		ram_buffer(14418) := X"00000000";
		ram_buffer(14419) := X"00000000";
		ram_buffer(14420) := X"00000000";
		ram_buffer(14421) := X"00000000";
		ram_buffer(14422) := X"00000000";
		ram_buffer(14423) := X"00000000";
		ram_buffer(14424) := X"00000000";
		ram_buffer(14425) := X"00000000";
		ram_buffer(14426) := X"00000000";
		ram_buffer(14427) := X"00000000";
		ram_buffer(14428) := X"00000000";
		ram_buffer(14429) := X"00000000";
		ram_buffer(14430) := X"00000000";
		ram_buffer(14431) := X"00000000";
		ram_buffer(14432) := X"00000000";
		ram_buffer(14433) := X"00000000";
		ram_buffer(14434) := X"00000000";
		ram_buffer(14435) := X"00000000";
		ram_buffer(14436) := X"00000000";
		ram_buffer(14437) := X"00000000";
		ram_buffer(14438) := X"00000000";
		ram_buffer(14439) := X"00000000";
		ram_buffer(14440) := X"00000000";
		ram_buffer(14441) := X"00000000";
		ram_buffer(14442) := X"00000000";
		ram_buffer(14443) := X"00000000";
		ram_buffer(14444) := X"00000000";
		ram_buffer(14445) := X"00000000";
		ram_buffer(14446) := X"00000000";
		ram_buffer(14447) := X"00000000";
		ram_buffer(14448) := X"00000000";
		ram_buffer(14449) := X"00000000";
		ram_buffer(14450) := X"00000000";
		ram_buffer(14451) := X"00000000";
		ram_buffer(14452) := X"00000000";
		ram_buffer(14453) := X"00000000";
		ram_buffer(14454) := X"00000000";
		ram_buffer(14455) := X"00000000";
		ram_buffer(14456) := X"00000000";
		ram_buffer(14457) := X"00000000";
		ram_buffer(14458) := X"00000000";
		ram_buffer(14459) := X"00000000";
		ram_buffer(14460) := X"00000000";
		ram_buffer(14461) := X"00000000";
		ram_buffer(14462) := X"00000000";
		ram_buffer(14463) := X"00000000";
		ram_buffer(14464) := X"00000000";
		ram_buffer(14465) := X"00000000";
		ram_buffer(14466) := X"00000000";
		ram_buffer(14467) := X"00000000";
		ram_buffer(14468) := X"00000000";
		ram_buffer(14469) := X"00000000";
		ram_buffer(14470) := X"00000000";
		ram_buffer(14471) := X"00000000";
		ram_buffer(14472) := X"00000000";
		ram_buffer(14473) := X"00000000";
		ram_buffer(14474) := X"00000000";
		ram_buffer(14475) := X"00000000";
		ram_buffer(14476) := X"00000000";
		ram_buffer(14477) := X"00000000";
		ram_buffer(14478) := X"00000000";
		ram_buffer(14479) := X"00000000";
		ram_buffer(14480) := X"00000000";
		ram_buffer(14481) := X"00000000";
		ram_buffer(14482) := X"00000000";
		ram_buffer(14483) := X"00000000";
		ram_buffer(14484) := X"00000000";
		ram_buffer(14485) := X"00000000";
		ram_buffer(14486) := X"00000000";
		ram_buffer(14487) := X"00000000";
		ram_buffer(14488) := X"00000000";
		ram_buffer(14489) := X"00000000";
		ram_buffer(14490) := X"00000000";
		ram_buffer(14491) := X"00000000";
		ram_buffer(14492) := X"00000000";
		ram_buffer(14493) := X"00000000";
		ram_buffer(14494) := X"00000000";
		ram_buffer(14495) := X"00000000";
		ram_buffer(14496) := X"00000000";
		ram_buffer(14497) := X"00000000";
		ram_buffer(14498) := X"00000000";
		ram_buffer(14499) := X"00000000";
		ram_buffer(14500) := X"00000000";
		ram_buffer(14501) := X"00000000";
		ram_buffer(14502) := X"00000000";
		ram_buffer(14503) := X"00000000";
		ram_buffer(14504) := X"00000000";
		ram_buffer(14505) := X"00000000";
		ram_buffer(14506) := X"00000000";
		ram_buffer(14507) := X"00000000";
		ram_buffer(14508) := X"00000000";
		ram_buffer(14509) := X"00000000";
		ram_buffer(14510) := X"00000000";
		ram_buffer(14511) := X"00000000";
		ram_buffer(14512) := X"00000000";
		ram_buffer(14513) := X"00000000";
		ram_buffer(14514) := X"00000000";
		ram_buffer(14515) := X"00000000";
		ram_buffer(14516) := X"00000000";
		ram_buffer(14517) := X"00000000";
		ram_buffer(14518) := X"00000000";
		ram_buffer(14519) := X"00000000";
		ram_buffer(14520) := X"00000000";
		ram_buffer(14521) := X"00000000";
		ram_buffer(14522) := X"00000000";
		ram_buffer(14523) := X"00000000";
		ram_buffer(14524) := X"00000000";
		ram_buffer(14525) := X"00000000";
		ram_buffer(14526) := X"00000000";
		ram_buffer(14527) := X"00000000";
		ram_buffer(14528) := X"00000000";
		ram_buffer(14529) := X"00000000";
		ram_buffer(14530) := X"00000000";
		ram_buffer(14531) := X"00000000";
		ram_buffer(14532) := X"00000000";
		ram_buffer(14533) := X"00000000";
		ram_buffer(14534) := X"00000000";
		ram_buffer(14535) := X"00000000";
		ram_buffer(14536) := X"00000000";
		ram_buffer(14537) := X"00000000";
		ram_buffer(14538) := X"00000000";
		ram_buffer(14539) := X"00000000";
		ram_buffer(14540) := X"00000000";
		ram_buffer(14541) := X"00000000";
		ram_buffer(14542) := X"00000000";
		ram_buffer(14543) := X"00000000";
		ram_buffer(14544) := X"00000000";
		ram_buffer(14545) := X"00000000";
		ram_buffer(14546) := X"00000000";
		ram_buffer(14547) := X"00000000";
		ram_buffer(14548) := X"00000000";
		ram_buffer(14549) := X"00000000";
		ram_buffer(14550) := X"00000000";
		ram_buffer(14551) := X"00000000";
		ram_buffer(14552) := X"00000000";
		ram_buffer(14553) := X"00000000";
		ram_buffer(14554) := X"00000000";
		ram_buffer(14555) := X"00000000";
		ram_buffer(14556) := X"00000000";
		ram_buffer(14557) := X"00000000";
		ram_buffer(14558) := X"00000000";
		ram_buffer(14559) := X"00000000";
		ram_buffer(14560) := X"00000000";
		ram_buffer(14561) := X"00000000";
		ram_buffer(14562) := X"00000000";
		ram_buffer(14563) := X"00000000";
		ram_buffer(14564) := X"00000000";
		ram_buffer(14565) := X"00000000";
		ram_buffer(14566) := X"00000000";
		ram_buffer(14567) := X"00000000";
		ram_buffer(14568) := X"00000000";
		ram_buffer(14569) := X"00000000";
		ram_buffer(14570) := X"00000000";
		ram_buffer(14571) := X"00000000";
		ram_buffer(14572) := X"00000000";
		ram_buffer(14573) := X"00000000";
		ram_buffer(14574) := X"00000000";
		ram_buffer(14575) := X"00000000";
		ram_buffer(14576) := X"00000000";
		ram_buffer(14577) := X"00000000";
		ram_buffer(14578) := X"00000000";
		ram_buffer(14579) := X"00000000";
		ram_buffer(14580) := X"00000000";
		ram_buffer(14581) := X"00000000";
		ram_buffer(14582) := X"00000000";
		ram_buffer(14583) := X"00000000";
		ram_buffer(14584) := X"00000000";
		ram_buffer(14585) := X"00000000";
		ram_buffer(14586) := X"00000000";
		ram_buffer(14587) := X"00000000";
		ram_buffer(14588) := X"00000000";
		ram_buffer(14589) := X"00000000";
		ram_buffer(14590) := X"00000000";
		ram_buffer(14591) := X"00000000";
		ram_buffer(14592) := X"00000000";
		ram_buffer(14593) := X"00000000";
		ram_buffer(14594) := X"00000000";
		ram_buffer(14595) := X"00000000";
		ram_buffer(14596) := X"00000000";
		ram_buffer(14597) := X"00000000";
		ram_buffer(14598) := X"00000000";
		ram_buffer(14599) := X"00000000";
		ram_buffer(14600) := X"00000000";
		ram_buffer(14601) := X"00000000";
		ram_buffer(14602) := X"00000000";
		ram_buffer(14603) := X"00000000";
		ram_buffer(14604) := X"00000000";
		ram_buffer(14605) := X"00000000";
		ram_buffer(14606) := X"00000000";
		ram_buffer(14607) := X"00000000";
		ram_buffer(14608) := X"00000000";
		ram_buffer(14609) := X"00000000";
		ram_buffer(14610) := X"00000000";
		ram_buffer(14611) := X"00000000";
		ram_buffer(14612) := X"00000000";
		ram_buffer(14613) := X"00000000";
		ram_buffer(14614) := X"00000000";
		ram_buffer(14615) := X"00000000";
		ram_buffer(14616) := X"00000000";
		ram_buffer(14617) := X"00000000";
		ram_buffer(14618) := X"00000000";
		ram_buffer(14619) := X"00000000";
		ram_buffer(14620) := X"00000000";
		ram_buffer(14621) := X"00000000";
		ram_buffer(14622) := X"00000000";
		ram_buffer(14623) := X"00000000";
		ram_buffer(14624) := X"00000000";
		ram_buffer(14625) := X"00000000";
		ram_buffer(14626) := X"00000000";
		ram_buffer(14627) := X"00000000";
		ram_buffer(14628) := X"00000000";
		ram_buffer(14629) := X"00000000";
		ram_buffer(14630) := X"00000000";
		ram_buffer(14631) := X"00000000";
		ram_buffer(14632) := X"00000000";
		ram_buffer(14633) := X"00000000";
		ram_buffer(14634) := X"00000000";
		ram_buffer(14635) := X"00000000";
		ram_buffer(14636) := X"00000000";
		ram_buffer(14637) := X"00000000";
		ram_buffer(14638) := X"00000000";
		ram_buffer(14639) := X"00000000";
		ram_buffer(14640) := X"00000000";
		ram_buffer(14641) := X"00000000";
		ram_buffer(14642) := X"00000000";
		ram_buffer(14643) := X"00000000";
		ram_buffer(14644) := X"00000000";
		ram_buffer(14645) := X"00000000";
		ram_buffer(14646) := X"00000000";
		ram_buffer(14647) := X"00000000";
		ram_buffer(14648) := X"00000000";
		ram_buffer(14649) := X"00000000";
		ram_buffer(14650) := X"00000000";
		ram_buffer(14651) := X"00000000";
		ram_buffer(14652) := X"00000000";
		ram_buffer(14653) := X"00000000";
		ram_buffer(14654) := X"00000000";
		ram_buffer(14655) := X"00000000";
		ram_buffer(14656) := X"00000000";
		ram_buffer(14657) := X"00000000";
		ram_buffer(14658) := X"00000000";
		ram_buffer(14659) := X"00000000";
		ram_buffer(14660) := X"00000000";
		ram_buffer(14661) := X"00000000";
		ram_buffer(14662) := X"00000000";
		ram_buffer(14663) := X"00000000";
		ram_buffer(14664) := X"00000000";
		ram_buffer(14665) := X"00000000";
		ram_buffer(14666) := X"00000000";
		ram_buffer(14667) := X"00000000";
		ram_buffer(14668) := X"00000000";
		ram_buffer(14669) := X"00000000";
		ram_buffer(14670) := X"00000000";
		ram_buffer(14671) := X"00000000";
		ram_buffer(14672) := X"00000000";
		ram_buffer(14673) := X"00000000";
		ram_buffer(14674) := X"00000000";
		ram_buffer(14675) := X"00000000";
		ram_buffer(14676) := X"00000000";
		ram_buffer(14677) := X"00000000";
		ram_buffer(14678) := X"00000000";
		ram_buffer(14679) := X"00000000";
		ram_buffer(14680) := X"00000000";
		ram_buffer(14681) := X"00000000";
		ram_buffer(14682) := X"00000000";
		ram_buffer(14683) := X"00000000";
		ram_buffer(14684) := X"00000000";
		ram_buffer(14685) := X"00000000";
		ram_buffer(14686) := X"00000000";
		ram_buffer(14687) := X"00000000";
		ram_buffer(14688) := X"00000000";
		ram_buffer(14689) := X"00000000";
		ram_buffer(14690) := X"00000000";
		ram_buffer(14691) := X"00000000";
		ram_buffer(14692) := X"00000000";
		ram_buffer(14693) := X"00000000";
		ram_buffer(14694) := X"00000000";
		ram_buffer(14695) := X"00000000";
		ram_buffer(14696) := X"00000000";
		ram_buffer(14697) := X"00000000";
		ram_buffer(14698) := X"00000000";
		ram_buffer(14699) := X"00000000";
		ram_buffer(14700) := X"00000000";
		ram_buffer(14701) := X"00000000";
		ram_buffer(14702) := X"00000000";
		ram_buffer(14703) := X"00000000";
		ram_buffer(14704) := X"00000000";
		ram_buffer(14705) := X"00000000";
		ram_buffer(14706) := X"00000000";
		ram_buffer(14707) := X"00000000";
		ram_buffer(14708) := X"00000000";
		ram_buffer(14709) := X"00000000";
		ram_buffer(14710) := X"00000000";
		ram_buffer(14711) := X"00000000";
		ram_buffer(14712) := X"00000000";
		ram_buffer(14713) := X"00000000";
		ram_buffer(14714) := X"00000000";
		ram_buffer(14715) := X"00000000";
		ram_buffer(14716) := X"00000000";
		ram_buffer(14717) := X"00000000";
		ram_buffer(14718) := X"00000000";
		ram_buffer(14719) := X"00000000";
		ram_buffer(14720) := X"00000000";
		ram_buffer(14721) := X"00000000";
		ram_buffer(14722) := X"00000000";
		ram_buffer(14723) := X"00000000";
		ram_buffer(14724) := X"00000000";
		ram_buffer(14725) := X"00000000";
		ram_buffer(14726) := X"00000000";
		ram_buffer(14727) := X"00000000";
		ram_buffer(14728) := X"00000000";
		ram_buffer(14729) := X"00000000";
		ram_buffer(14730) := X"00000000";
		ram_buffer(14731) := X"00000000";
		ram_buffer(14732) := X"00000000";
		ram_buffer(14733) := X"00000000";
		ram_buffer(14734) := X"00000000";
		ram_buffer(14735) := X"00000000";
		ram_buffer(14736) := X"00000000";
		ram_buffer(14737) := X"00000000";
		ram_buffer(14738) := X"00000000";
		ram_buffer(14739) := X"00000000";
		ram_buffer(14740) := X"00000000";
		ram_buffer(14741) := X"00000000";
		ram_buffer(14742) := X"00000000";
		ram_buffer(14743) := X"00000000";
		ram_buffer(14744) := X"00000000";
		ram_buffer(14745) := X"00000000";
		ram_buffer(14746) := X"00000000";
		ram_buffer(14747) := X"00000000";
		ram_buffer(14748) := X"00000000";
		ram_buffer(14749) := X"00000000";
		ram_buffer(14750) := X"00000000";
		ram_buffer(14751) := X"00000000";
		ram_buffer(14752) := X"00000000";
		ram_buffer(14753) := X"00000000";
		ram_buffer(14754) := X"00000000";
		ram_buffer(14755) := X"00000000";
		ram_buffer(14756) := X"00000000";
		ram_buffer(14757) := X"00000000";
		ram_buffer(14758) := X"00000000";
		ram_buffer(14759) := X"00000000";
		ram_buffer(14760) := X"00000000";
		ram_buffer(14761) := X"00000000";
		ram_buffer(14762) := X"00000000";
		ram_buffer(14763) := X"00000000";
		ram_buffer(14764) := X"00000000";
		ram_buffer(14765) := X"00000000";
		ram_buffer(14766) := X"00000000";
		ram_buffer(14767) := X"00000000";
		ram_buffer(14768) := X"00000000";
		ram_buffer(14769) := X"00000000";
		ram_buffer(14770) := X"00000000";
		ram_buffer(14771) := X"00000000";
		ram_buffer(14772) := X"00000000";
		ram_buffer(14773) := X"00000000";
		ram_buffer(14774) := X"00000000";
		ram_buffer(14775) := X"00000000";
		ram_buffer(14776) := X"00000000";
		ram_buffer(14777) := X"00000000";
		ram_buffer(14778) := X"00000000";
		ram_buffer(14779) := X"00000000";
		ram_buffer(14780) := X"00000000";
		ram_buffer(14781) := X"00000000";
		ram_buffer(14782) := X"00000000";
		ram_buffer(14783) := X"00000000";
		ram_buffer(14784) := X"00000000";
		ram_buffer(14785) := X"00000000";
		ram_buffer(14786) := X"00000000";
		ram_buffer(14787) := X"00000000";
		ram_buffer(14788) := X"00000000";
		ram_buffer(14789) := X"00000000";
		ram_buffer(14790) := X"00000000";
		ram_buffer(14791) := X"00000000";
		ram_buffer(14792) := X"00000000";
		ram_buffer(14793) := X"00000000";
		ram_buffer(14794) := X"00000000";
		ram_buffer(14795) := X"00000000";
		ram_buffer(14796) := X"00000000";
		ram_buffer(14797) := X"00000000";
		ram_buffer(14798) := X"00000000";
		ram_buffer(14799) := X"00000000";
		ram_buffer(14800) := X"00000000";
		ram_buffer(14801) := X"00000000";
		ram_buffer(14802) := X"00000000";
		ram_buffer(14803) := X"00000000";
		ram_buffer(14804) := X"00000000";
		ram_buffer(14805) := X"00000000";
		ram_buffer(14806) := X"00000000";
		ram_buffer(14807) := X"00000000";
		ram_buffer(14808) := X"00000000";
		ram_buffer(14809) := X"00000000";
		ram_buffer(14810) := X"00000000";
		ram_buffer(14811) := X"00000000";
		ram_buffer(14812) := X"00000000";
		ram_buffer(14813) := X"00000000";
		ram_buffer(14814) := X"00000000";
		ram_buffer(14815) := X"00000000";
		ram_buffer(14816) := X"00000000";
		ram_buffer(14817) := X"00000000";
		ram_buffer(14818) := X"00000000";
		ram_buffer(14819) := X"00000000";
		ram_buffer(14820) := X"00000000";
		ram_buffer(14821) := X"00000000";
		ram_buffer(14822) := X"00000000";
		ram_buffer(14823) := X"00000000";
		ram_buffer(14824) := X"00000000";
		ram_buffer(14825) := X"00000000";
		ram_buffer(14826) := X"00000000";
		ram_buffer(14827) := X"00000000";
		ram_buffer(14828) := X"00000000";
		ram_buffer(14829) := X"00000000";
		ram_buffer(14830) := X"00000000";
		ram_buffer(14831) := X"00000000";
		ram_buffer(14832) := X"00000000";
		ram_buffer(14833) := X"00000000";
		ram_buffer(14834) := X"00000000";
		ram_buffer(14835) := X"00000000";
		ram_buffer(14836) := X"00000000";
		ram_buffer(14837) := X"00000000";
		ram_buffer(14838) := X"00000000";
		ram_buffer(14839) := X"00000000";
		ram_buffer(14840) := X"00000000";
		ram_buffer(14841) := X"00000000";
		ram_buffer(14842) := X"00000000";
		ram_buffer(14843) := X"00000000";
		ram_buffer(14844) := X"00000000";
		ram_buffer(14845) := X"00000000";
		ram_buffer(14846) := X"00000000";
		ram_buffer(14847) := X"00000000";
		ram_buffer(14848) := X"00000000";
		ram_buffer(14849) := X"00000000";
		ram_buffer(14850) := X"00000000";
		ram_buffer(14851) := X"00000000";
		ram_buffer(14852) := X"00000000";
		ram_buffer(14853) := X"00000000";
		ram_buffer(14854) := X"00000000";
		ram_buffer(14855) := X"00000000";
		ram_buffer(14856) := X"00000000";
		ram_buffer(14857) := X"00000000";
		ram_buffer(14858) := X"00000000";
		ram_buffer(14859) := X"00000000";
		ram_buffer(14860) := X"00000000";
		ram_buffer(14861) := X"00000000";
		ram_buffer(14862) := X"00000000";
		ram_buffer(14863) := X"00000000";
		ram_buffer(14864) := X"00000000";
		ram_buffer(14865) := X"00000000";
		ram_buffer(14866) := X"00000000";
		ram_buffer(14867) := X"00000000";
		ram_buffer(14868) := X"00000000";
		ram_buffer(14869) := X"00000000";
		ram_buffer(14870) := X"00000000";
		ram_buffer(14871) := X"00000000";
		ram_buffer(14872) := X"00000000";
		ram_buffer(14873) := X"00000000";
		ram_buffer(14874) := X"00000000";
		ram_buffer(14875) := X"00000000";
		ram_buffer(14876) := X"00000000";
		ram_buffer(14877) := X"00000000";
		ram_buffer(14878) := X"00000000";
		ram_buffer(14879) := X"00000000";
		ram_buffer(14880) := X"00000000";
		ram_buffer(14881) := X"00000000";
		ram_buffer(14882) := X"00000000";
		ram_buffer(14883) := X"00000000";
		ram_buffer(14884) := X"00000000";
		ram_buffer(14885) := X"00000000";
		ram_buffer(14886) := X"00000000";
		ram_buffer(14887) := X"00000000";
		ram_buffer(14888) := X"00000000";
		ram_buffer(14889) := X"00000000";
		ram_buffer(14890) := X"00000000";
		ram_buffer(14891) := X"00000000";
		ram_buffer(14892) := X"00000000";
		ram_buffer(14893) := X"00000000";
		ram_buffer(14894) := X"00000000";
		ram_buffer(14895) := X"00000000";
		ram_buffer(14896) := X"00000000";
		ram_buffer(14897) := X"00000000";
		ram_buffer(14898) := X"00000000";
		ram_buffer(14899) := X"00000000";
		ram_buffer(14900) := X"00000000";
		ram_buffer(14901) := X"00000000";
		ram_buffer(14902) := X"00000000";
		ram_buffer(14903) := X"00000000";
		ram_buffer(14904) := X"00000000";
		ram_buffer(14905) := X"00000000";
		ram_buffer(14906) := X"00000000";
		ram_buffer(14907) := X"00000000";
		ram_buffer(14908) := X"00000000";
		ram_buffer(14909) := X"00000000";
		ram_buffer(14910) := X"00000000";
		ram_buffer(14911) := X"00000000";
		ram_buffer(14912) := X"00000000";
		ram_buffer(14913) := X"00000000";
		ram_buffer(14914) := X"00000000";
		ram_buffer(14915) := X"00000000";
		ram_buffer(14916) := X"00000000";
		ram_buffer(14917) := X"00000000";
		ram_buffer(14918) := X"00000000";
		ram_buffer(14919) := X"00000000";
		ram_buffer(14920) := X"00000000";
		ram_buffer(14921) := X"00000000";
		ram_buffer(14922) := X"00000000";
		ram_buffer(14923) := X"00000000";
		ram_buffer(14924) := X"00000000";
		ram_buffer(14925) := X"00000000";
		ram_buffer(14926) := X"00000000";
		ram_buffer(14927) := X"00000000";
		ram_buffer(14928) := X"00000000";
		ram_buffer(14929) := X"00000000";
		ram_buffer(14930) := X"00000000";
		ram_buffer(14931) := X"00000000";
		ram_buffer(14932) := X"00000000";
		ram_buffer(14933) := X"00000000";
		ram_buffer(14934) := X"00000000";
		ram_buffer(14935) := X"00000000";
		ram_buffer(14936) := X"00000000";
		ram_buffer(14937) := X"00000000";
		ram_buffer(14938) := X"00000000";
		ram_buffer(14939) := X"00000000";
		ram_buffer(14940) := X"00000000";
		ram_buffer(14941) := X"00000000";
		ram_buffer(14942) := X"00000000";
		ram_buffer(14943) := X"00000000";
		ram_buffer(14944) := X"00000000";
		ram_buffer(14945) := X"00000000";
		ram_buffer(14946) := X"00000000";
		ram_buffer(14947) := X"00000000";
		ram_buffer(14948) := X"00000000";
		ram_buffer(14949) := X"00000000";
		ram_buffer(14950) := X"00000000";
		ram_buffer(14951) := X"00000000";
		ram_buffer(14952) := X"00000000";
		ram_buffer(14953) := X"00000000";
		ram_buffer(14954) := X"00000000";
		ram_buffer(14955) := X"00000000";
		ram_buffer(14956) := X"00000000";
		ram_buffer(14957) := X"00000000";
		ram_buffer(14958) := X"00000000";
		ram_buffer(14959) := X"00000000";
		ram_buffer(14960) := X"00000000";
		ram_buffer(14961) := X"00000000";
		ram_buffer(14962) := X"00000000";
		ram_buffer(14963) := X"00000000";
		ram_buffer(14964) := X"00000000";
		ram_buffer(14965) := X"00000000";
		ram_buffer(14966) := X"00000000";
		ram_buffer(14967) := X"00000000";
		ram_buffer(14968) := X"00000000";
		ram_buffer(14969) := X"00000000";
		ram_buffer(14970) := X"00000000";
		ram_buffer(14971) := X"00000000";
		ram_buffer(14972) := X"00000000";
		ram_buffer(14973) := X"00000000";
		ram_buffer(14974) := X"00000000";
		ram_buffer(14975) := X"00000000";
		ram_buffer(14976) := X"00000000";
		ram_buffer(14977) := X"00000000";
		ram_buffer(14978) := X"00000000";
		ram_buffer(14979) := X"00000000";
		ram_buffer(14980) := X"00000000";
		ram_buffer(14981) := X"00000000";
		ram_buffer(14982) := X"00000000";
		ram_buffer(14983) := X"00000000";
		ram_buffer(14984) := X"00000000";
		ram_buffer(14985) := X"00000000";
		ram_buffer(14986) := X"00000000";
		ram_buffer(14987) := X"00000000";
		ram_buffer(14988) := X"00000000";
		ram_buffer(14989) := X"00000000";
		ram_buffer(14990) := X"00000000";
		ram_buffer(14991) := X"00000000";
		ram_buffer(14992) := X"00000000";
		ram_buffer(14993) := X"00000000";
		ram_buffer(14994) := X"00000000";
		ram_buffer(14995) := X"00000000";
		ram_buffer(14996) := X"00000000";
		ram_buffer(14997) := X"00000000";
		ram_buffer(14998) := X"00000000";
		ram_buffer(14999) := X"00000000";
		ram_buffer(15000) := X"00000000";
		ram_buffer(15001) := X"00000000";
		ram_buffer(15002) := X"00000000";
		ram_buffer(15003) := X"00000000";
		ram_buffer(15004) := X"00000000";
		ram_buffer(15005) := X"00000000";
		ram_buffer(15006) := X"00000000";
		ram_buffer(15007) := X"00000000";
		ram_buffer(15008) := X"00000000";
		ram_buffer(15009) := X"00000000";
		ram_buffer(15010) := X"00000000";
		ram_buffer(15011) := X"00000000";
		ram_buffer(15012) := X"00000000";
		ram_buffer(15013) := X"00000000";
		ram_buffer(15014) := X"00000000";
		ram_buffer(15015) := X"00000000";
		ram_buffer(15016) := X"00000000";
		ram_buffer(15017) := X"00000000";
		ram_buffer(15018) := X"00000000";
		ram_buffer(15019) := X"00000000";
		ram_buffer(15020) := X"00000000";
		ram_buffer(15021) := X"00000000";
		ram_buffer(15022) := X"00000000";
		ram_buffer(15023) := X"00000000";
		ram_buffer(15024) := X"00000000";
		ram_buffer(15025) := X"00000000";
		ram_buffer(15026) := X"00000000";
		ram_buffer(15027) := X"00000000";
		ram_buffer(15028) := X"00000000";
		ram_buffer(15029) := X"00000000";
		ram_buffer(15030) := X"00000000";
		ram_buffer(15031) := X"00000000";
		ram_buffer(15032) := X"00000000";
		ram_buffer(15033) := X"00000000";
		ram_buffer(15034) := X"00000000";
		ram_buffer(15035) := X"00000000";
		ram_buffer(15036) := X"00000000";
		ram_buffer(15037) := X"00000000";
		ram_buffer(15038) := X"00000000";
		ram_buffer(15039) := X"00000000";
		ram_buffer(15040) := X"00000000";
		ram_buffer(15041) := X"00000000";
		ram_buffer(15042) := X"00000000";
		ram_buffer(15043) := X"00000000";
		ram_buffer(15044) := X"00000000";
		ram_buffer(15045) := X"00000000";
		ram_buffer(15046) := X"00000000";
		ram_buffer(15047) := X"00000000";
		ram_buffer(15048) := X"00000000";
		ram_buffer(15049) := X"00000000";
		ram_buffer(15050) := X"00000000";
		ram_buffer(15051) := X"00000000";
		ram_buffer(15052) := X"00000000";
		ram_buffer(15053) := X"00000000";
		ram_buffer(15054) := X"00000000";
		ram_buffer(15055) := X"00000000";
		ram_buffer(15056) := X"00000000";
		ram_buffer(15057) := X"00000000";
		ram_buffer(15058) := X"00000000";
		ram_buffer(15059) := X"00000000";
		ram_buffer(15060) := X"00000000";
		ram_buffer(15061) := X"00000000";
		ram_buffer(15062) := X"00000000";
		ram_buffer(15063) := X"00000000";
		ram_buffer(15064) := X"00000000";
		ram_buffer(15065) := X"00000000";
		ram_buffer(15066) := X"00000000";
		ram_buffer(15067) := X"00000000";
		ram_buffer(15068) := X"00000000";
		ram_buffer(15069) := X"00000000";
		ram_buffer(15070) := X"00000000";
		ram_buffer(15071) := X"00000000";
		ram_buffer(15072) := X"00000000";
		ram_buffer(15073) := X"00000000";
		ram_buffer(15074) := X"00000000";
		ram_buffer(15075) := X"00000000";
		ram_buffer(15076) := X"00000000";
		ram_buffer(15077) := X"00000000";
		ram_buffer(15078) := X"00000000";
		ram_buffer(15079) := X"00000000";
		ram_buffer(15080) := X"00000000";
		ram_buffer(15081) := X"00000000";
		ram_buffer(15082) := X"00000000";
		ram_buffer(15083) := X"00000000";
		ram_buffer(15084) := X"00000000";
		ram_buffer(15085) := X"00000000";
		ram_buffer(15086) := X"00000000";
		ram_buffer(15087) := X"00000000";
		ram_buffer(15088) := X"00000000";
		ram_buffer(15089) := X"00000000";
		ram_buffer(15090) := X"00000000";
		ram_buffer(15091) := X"00000000";
		ram_buffer(15092) := X"00000000";
		ram_buffer(15093) := X"00000000";
		ram_buffer(15094) := X"00000000";
		ram_buffer(15095) := X"00000000";
		ram_buffer(15096) := X"00000000";
		ram_buffer(15097) := X"00000000";
		ram_buffer(15098) := X"00000000";
		ram_buffer(15099) := X"00000000";
		ram_buffer(15100) := X"00000000";
		ram_buffer(15101) := X"00000000";
		ram_buffer(15102) := X"00000000";
		ram_buffer(15103) := X"00000000";
		ram_buffer(15104) := X"00000000";
		ram_buffer(15105) := X"00000000";
		ram_buffer(15106) := X"00000000";
		ram_buffer(15107) := X"00000000";
		ram_buffer(15108) := X"00000000";
		ram_buffer(15109) := X"00000000";
		ram_buffer(15110) := X"00000000";
		ram_buffer(15111) := X"00000000";
		ram_buffer(15112) := X"00000000";
		ram_buffer(15113) := X"00000000";
		ram_buffer(15114) := X"00000000";
		ram_buffer(15115) := X"00000000";
		ram_buffer(15116) := X"00000000";
		ram_buffer(15117) := X"00000000";
		ram_buffer(15118) := X"00000000";
		ram_buffer(15119) := X"00000000";
		ram_buffer(15120) := X"00000000";
		ram_buffer(15121) := X"00000000";
		ram_buffer(15122) := X"00000000";
		ram_buffer(15123) := X"00000000";
		ram_buffer(15124) := X"00000000";
		ram_buffer(15125) := X"00000000";
		ram_buffer(15126) := X"00000000";
		ram_buffer(15127) := X"00000000";
		ram_buffer(15128) := X"00000000";
		ram_buffer(15129) := X"00000000";
		ram_buffer(15130) := X"00000000";
		ram_buffer(15131) := X"00000000";
		ram_buffer(15132) := X"00000000";
		ram_buffer(15133) := X"00000000";
		ram_buffer(15134) := X"00000000";
		ram_buffer(15135) := X"00000000";
		ram_buffer(15136) := X"00000000";
		ram_buffer(15137) := X"00000000";
		ram_buffer(15138) := X"00000000";
		ram_buffer(15139) := X"00000000";
		ram_buffer(15140) := X"00000000";
		ram_buffer(15141) := X"00000000";
		ram_buffer(15142) := X"00000000";
		ram_buffer(15143) := X"00000000";
		ram_buffer(15144) := X"00000000";
		ram_buffer(15145) := X"00000000";
		ram_buffer(15146) := X"00000000";
		ram_buffer(15147) := X"00000000";
		ram_buffer(15148) := X"00000000";
		ram_buffer(15149) := X"00000000";
		ram_buffer(15150) := X"00000000";
		ram_buffer(15151) := X"00000000";
		ram_buffer(15152) := X"00000000";
		ram_buffer(15153) := X"00000000";
		ram_buffer(15154) := X"00000000";
		ram_buffer(15155) := X"00000000";
		ram_buffer(15156) := X"00000000";
		ram_buffer(15157) := X"00000000";
		ram_buffer(15158) := X"00000000";
		ram_buffer(15159) := X"00000000";
		ram_buffer(15160) := X"00000000";
		ram_buffer(15161) := X"00000000";
		ram_buffer(15162) := X"00000000";
		ram_buffer(15163) := X"00000000";
		ram_buffer(15164) := X"00000000";
		ram_buffer(15165) := X"00000000";
		ram_buffer(15166) := X"00000000";
		ram_buffer(15167) := X"00000000";
		ram_buffer(15168) := X"00000000";
		ram_buffer(15169) := X"00000000";
		ram_buffer(15170) := X"00000000";
		ram_buffer(15171) := X"00000000";
		ram_buffer(15172) := X"00000000";
		ram_buffer(15173) := X"00000000";
		ram_buffer(15174) := X"00000000";
		ram_buffer(15175) := X"00000000";
		ram_buffer(15176) := X"00000000";
		ram_buffer(15177) := X"00000000";
		ram_buffer(15178) := X"00000000";
		ram_buffer(15179) := X"00000000";
		ram_buffer(15180) := X"00000000";
		ram_buffer(15181) := X"00000000";
		ram_buffer(15182) := X"00000000";
		ram_buffer(15183) := X"00000000";
		ram_buffer(15184) := X"00000000";
		ram_buffer(15185) := X"00000000";
		ram_buffer(15186) := X"00000000";
		ram_buffer(15187) := X"00000000";
		ram_buffer(15188) := X"00000000";
		ram_buffer(15189) := X"00000000";
		ram_buffer(15190) := X"00000000";
		ram_buffer(15191) := X"00000000";
		ram_buffer(15192) := X"00000000";
		ram_buffer(15193) := X"00000000";
		ram_buffer(15194) := X"00000000";
		ram_buffer(15195) := X"00000000";
		ram_buffer(15196) := X"00000000";
		ram_buffer(15197) := X"00000000";
		ram_buffer(15198) := X"00000000";
		ram_buffer(15199) := X"00000000";
		ram_buffer(15200) := X"00000000";
		ram_buffer(15201) := X"00000000";
		ram_buffer(15202) := X"00000000";
		ram_buffer(15203) := X"00000000";
		ram_buffer(15204) := X"00000000";
		ram_buffer(15205) := X"00000000";
		ram_buffer(15206) := X"00000000";
		ram_buffer(15207) := X"00000000";
		ram_buffer(15208) := X"00000000";
		ram_buffer(15209) := X"00000000";
		ram_buffer(15210) := X"00000000";
		ram_buffer(15211) := X"00000000";
		ram_buffer(15212) := X"00000000";
		ram_buffer(15213) := X"00000000";
		ram_buffer(15214) := X"00000000";
		ram_buffer(15215) := X"00000000";
		ram_buffer(15216) := X"00000000";
		ram_buffer(15217) := X"00000000";
		ram_buffer(15218) := X"00000000";
		ram_buffer(15219) := X"00000000";
		ram_buffer(15220) := X"00000000";
		ram_buffer(15221) := X"00000000";
		ram_buffer(15222) := X"00000000";
		ram_buffer(15223) := X"00000000";
		ram_buffer(15224) := X"00000000";
		ram_buffer(15225) := X"00000000";
		ram_buffer(15226) := X"00000000";
		ram_buffer(15227) := X"00000000";
		ram_buffer(15228) := X"00000000";
		ram_buffer(15229) := X"00000000";
		ram_buffer(15230) := X"00000000";
		ram_buffer(15231) := X"00000000";
		ram_buffer(15232) := X"00000000";
		ram_buffer(15233) := X"00000000";
		ram_buffer(15234) := X"00000000";
		ram_buffer(15235) := X"00000000";
		ram_buffer(15236) := X"00000000";
		ram_buffer(15237) := X"00000000";
		ram_buffer(15238) := X"00000000";
		ram_buffer(15239) := X"00000000";
		ram_buffer(15240) := X"00000000";
		ram_buffer(15241) := X"00000000";
		ram_buffer(15242) := X"00000000";
		ram_buffer(15243) := X"00000000";
		ram_buffer(15244) := X"00000000";
		ram_buffer(15245) := X"00000000";
		ram_buffer(15246) := X"00000000";
		ram_buffer(15247) := X"00000000";
		ram_buffer(15248) := X"00000000";
		ram_buffer(15249) := X"00000000";
		ram_buffer(15250) := X"00000000";
		ram_buffer(15251) := X"00000000";
		ram_buffer(15252) := X"00000000";
		ram_buffer(15253) := X"00000000";
		ram_buffer(15254) := X"00000000";
		ram_buffer(15255) := X"00000000";
		ram_buffer(15256) := X"00000000";
		ram_buffer(15257) := X"00000000";
		ram_buffer(15258) := X"00000000";
		ram_buffer(15259) := X"00000000";
		ram_buffer(15260) := X"00000000";
		ram_buffer(15261) := X"00000000";
		ram_buffer(15262) := X"00000000";
		ram_buffer(15263) := X"00000000";
		ram_buffer(15264) := X"00000000";
		ram_buffer(15265) := X"00000000";
		ram_buffer(15266) := X"00000000";
		ram_buffer(15267) := X"00000000";
		ram_buffer(15268) := X"00000000";
		ram_buffer(15269) := X"00000000";
		ram_buffer(15270) := X"00000000";
		ram_buffer(15271) := X"00000000";
		ram_buffer(15272) := X"00000000";
		ram_buffer(15273) := X"00000000";
		ram_buffer(15274) := X"00000000";
		ram_buffer(15275) := X"00000000";
		ram_buffer(15276) := X"00000000";
		ram_buffer(15277) := X"00000000";
		ram_buffer(15278) := X"00000000";
		ram_buffer(15279) := X"00000000";
		ram_buffer(15280) := X"00000000";
		ram_buffer(15281) := X"00000000";
		ram_buffer(15282) := X"00000000";
		ram_buffer(15283) := X"00000000";
		ram_buffer(15284) := X"00000000";
		ram_buffer(15285) := X"00000000";
		ram_buffer(15286) := X"00000000";
		ram_buffer(15287) := X"00000000";
		ram_buffer(15288) := X"00000000";
		ram_buffer(15289) := X"00000000";
		ram_buffer(15290) := X"00000000";
		ram_buffer(15291) := X"00000000";
		ram_buffer(15292) := X"00000000";
		ram_buffer(15293) := X"00000000";
		ram_buffer(15294) := X"00000000";
		ram_buffer(15295) := X"00000000";
		ram_buffer(15296) := X"00000000";
		ram_buffer(15297) := X"00000000";
		ram_buffer(15298) := X"00000000";
		ram_buffer(15299) := X"00000000";
		ram_buffer(15300) := X"00000000";
		ram_buffer(15301) := X"00000000";
		ram_buffer(15302) := X"00000000";
		ram_buffer(15303) := X"00000000";
		ram_buffer(15304) := X"00000000";
		ram_buffer(15305) := X"00000000";
		ram_buffer(15306) := X"00000000";
		ram_buffer(15307) := X"00000000";
		ram_buffer(15308) := X"00000000";
		ram_buffer(15309) := X"00000000";
		ram_buffer(15310) := X"00000000";
		ram_buffer(15311) := X"00000000";
		ram_buffer(15312) := X"00000000";
		ram_buffer(15313) := X"00000000";
		ram_buffer(15314) := X"00000000";
		ram_buffer(15315) := X"00000000";
		ram_buffer(15316) := X"00000000";
		ram_buffer(15317) := X"00000000";
		ram_buffer(15318) := X"00000000";
		ram_buffer(15319) := X"00000000";
		ram_buffer(15320) := X"00000000";
		ram_buffer(15321) := X"00000000";
		ram_buffer(15322) := X"00000000";
		ram_buffer(15323) := X"00000000";
		ram_buffer(15324) := X"00000000";
		ram_buffer(15325) := X"00000000";
		ram_buffer(15326) := X"00000000";
		ram_buffer(15327) := X"00000000";
		ram_buffer(15328) := X"00000000";
		ram_buffer(15329) := X"00000000";
		ram_buffer(15330) := X"00000000";
		ram_buffer(15331) := X"00000000";
		ram_buffer(15332) := X"00000000";
		ram_buffer(15333) := X"00000000";
		ram_buffer(15334) := X"00000000";
		ram_buffer(15335) := X"00000000";
		ram_buffer(15336) := X"00000000";
		ram_buffer(15337) := X"00000000";
		ram_buffer(15338) := X"00000000";
		ram_buffer(15339) := X"00000000";
		ram_buffer(15340) := X"00000000";
		ram_buffer(15341) := X"00000000";
		ram_buffer(15342) := X"00000000";
		ram_buffer(15343) := X"00000000";
		ram_buffer(15344) := X"00000000";
		ram_buffer(15345) := X"00000000";
		ram_buffer(15346) := X"00000000";
		ram_buffer(15347) := X"00000000";
		ram_buffer(15348) := X"00000000";
		ram_buffer(15349) := X"00000000";
		ram_buffer(15350) := X"00000000";
		ram_buffer(15351) := X"00000000";
		ram_buffer(15352) := X"00000000";
		ram_buffer(15353) := X"00000000";
		ram_buffer(15354) := X"00000000";
		ram_buffer(15355) := X"00000000";
		ram_buffer(15356) := X"00000000";
		ram_buffer(15357) := X"00000000";
		ram_buffer(15358) := X"00000000";
		ram_buffer(15359) := X"00000000";
		ram_buffer(15360) := X"00000000";
		ram_buffer(15361) := X"00000000";
		ram_buffer(15362) := X"00000000";
		ram_buffer(15363) := X"00000000";
		ram_buffer(15364) := X"00000000";
		ram_buffer(15365) := X"00000000";
		ram_buffer(15366) := X"00000000";
		ram_buffer(15367) := X"00000000";
		ram_buffer(15368) := X"00000000";
		ram_buffer(15369) := X"00000000";
		ram_buffer(15370) := X"00000000";
		ram_buffer(15371) := X"00000000";
		ram_buffer(15372) := X"00000000";
		ram_buffer(15373) := X"00000000";
		ram_buffer(15374) := X"00000000";
		ram_buffer(15375) := X"00000000";
		ram_buffer(15376) := X"00000000";
		ram_buffer(15377) := X"00000000";
		ram_buffer(15378) := X"00000000";
		ram_buffer(15379) := X"00000000";
		ram_buffer(15380) := X"00000000";
		ram_buffer(15381) := X"00000000";
		ram_buffer(15382) := X"00000000";
		ram_buffer(15383) := X"00000000";
		ram_buffer(15384) := X"00000000";
		ram_buffer(15385) := X"00000000";
		ram_buffer(15386) := X"00000000";
		ram_buffer(15387) := X"00000000";
		ram_buffer(15388) := X"00000000";
		ram_buffer(15389) := X"00000000";
		ram_buffer(15390) := X"00000000";
		ram_buffer(15391) := X"00000000";
		ram_buffer(15392) := X"00000000";
		ram_buffer(15393) := X"00000000";
		ram_buffer(15394) := X"00000000";
		ram_buffer(15395) := X"00000000";
		ram_buffer(15396) := X"00000000";
		ram_buffer(15397) := X"00000000";
		ram_buffer(15398) := X"00000000";
		ram_buffer(15399) := X"00000000";
		ram_buffer(15400) := X"00000000";
		ram_buffer(15401) := X"00000000";
		ram_buffer(15402) := X"00000000";
		ram_buffer(15403) := X"00000000";
		ram_buffer(15404) := X"00000000";
		ram_buffer(15405) := X"00000000";
		ram_buffer(15406) := X"00000000";
		ram_buffer(15407) := X"00000000";
		ram_buffer(15408) := X"00000000";
		ram_buffer(15409) := X"00000000";
		ram_buffer(15410) := X"00000000";
		ram_buffer(15411) := X"00000000";
		ram_buffer(15412) := X"00000000";
		ram_buffer(15413) := X"00000000";
		ram_buffer(15414) := X"00000000";
		ram_buffer(15415) := X"00000000";
		ram_buffer(15416) := X"00000000";
		ram_buffer(15417) := X"00000000";
		ram_buffer(15418) := X"00000000";
		ram_buffer(15419) := X"00000000";
		ram_buffer(15420) := X"00000000";
		ram_buffer(15421) := X"00000000";
		ram_buffer(15422) := X"00000000";
		ram_buffer(15423) := X"00000000";
		ram_buffer(15424) := X"00000000";
		ram_buffer(15425) := X"00000000";
		ram_buffer(15426) := X"00000000";
		ram_buffer(15427) := X"00000000";
		ram_buffer(15428) := X"00000000";
		ram_buffer(15429) := X"00000000";
		ram_buffer(15430) := X"00000000";
		ram_buffer(15431) := X"00000000";
		ram_buffer(15432) := X"00000000";
		ram_buffer(15433) := X"00000000";
		ram_buffer(15434) := X"00000000";
		ram_buffer(15435) := X"00000000";
		ram_buffer(15436) := X"00000000";
		ram_buffer(15437) := X"00000000";
		ram_buffer(15438) := X"00000000";
		ram_buffer(15439) := X"00000000";
		ram_buffer(15440) := X"00000000";
		ram_buffer(15441) := X"00000000";
		ram_buffer(15442) := X"00000000";
		ram_buffer(15443) := X"00000000";
		ram_buffer(15444) := X"00000000";
		ram_buffer(15445) := X"00000000";
		ram_buffer(15446) := X"00000000";
		ram_buffer(15447) := X"00000000";
		ram_buffer(15448) := X"00000000";
		ram_buffer(15449) := X"00000000";
		ram_buffer(15450) := X"00000000";
		ram_buffer(15451) := X"00000000";
		ram_buffer(15452) := X"00000000";
		ram_buffer(15453) := X"00000000";
		ram_buffer(15454) := X"00000000";
		ram_buffer(15455) := X"00000000";
		ram_buffer(15456) := X"00000000";
		ram_buffer(15457) := X"00000000";
		ram_buffer(15458) := X"00000000";
		ram_buffer(15459) := X"00000000";
		ram_buffer(15460) := X"00000000";
		ram_buffer(15461) := X"00000000";
		ram_buffer(15462) := X"00000000";
		ram_buffer(15463) := X"00000000";
		ram_buffer(15464) := X"00000000";
		ram_buffer(15465) := X"00000000";
		ram_buffer(15466) := X"00000000";
		ram_buffer(15467) := X"00000000";
		ram_buffer(15468) := X"00000000";
		ram_buffer(15469) := X"00000000";
		ram_buffer(15470) := X"00000000";
		ram_buffer(15471) := X"00000000";
		ram_buffer(15472) := X"00000000";
		ram_buffer(15473) := X"00000000";
		ram_buffer(15474) := X"00000000";
		ram_buffer(15475) := X"00000000";
		ram_buffer(15476) := X"00000000";
		ram_buffer(15477) := X"00000000";
		ram_buffer(15478) := X"00000000";
		ram_buffer(15479) := X"00000000";
		ram_buffer(15480) := X"00000000";
		ram_buffer(15481) := X"00000000";
		ram_buffer(15482) := X"00000000";
		ram_buffer(15483) := X"00000000";
		ram_buffer(15484) := X"00000000";
		ram_buffer(15485) := X"00000000";
		ram_buffer(15486) := X"00000000";
		ram_buffer(15487) := X"00000000";
		ram_buffer(15488) := X"00000000";
		ram_buffer(15489) := X"00000000";
		ram_buffer(15490) := X"00000000";
		ram_buffer(15491) := X"00000000";
		ram_buffer(15492) := X"00000000";
		ram_buffer(15493) := X"00000000";
		ram_buffer(15494) := X"00000000";
		ram_buffer(15495) := X"00000000";
		ram_buffer(15496) := X"00000000";
		ram_buffer(15497) := X"00000000";
		ram_buffer(15498) := X"00000000";
		ram_buffer(15499) := X"00000000";
		ram_buffer(15500) := X"00000000";
		ram_buffer(15501) := X"00000000";
		ram_buffer(15502) := X"00000000";
		ram_buffer(15503) := X"00000000";
		ram_buffer(15504) := X"00000000";
		ram_buffer(15505) := X"00000000";
		ram_buffer(15506) := X"00000000";
		ram_buffer(15507) := X"00000000";
		ram_buffer(15508) := X"00000000";
		ram_buffer(15509) := X"00000000";
		ram_buffer(15510) := X"00000000";
		ram_buffer(15511) := X"00000000";
		ram_buffer(15512) := X"00000000";
		ram_buffer(15513) := X"00000000";
		ram_buffer(15514) := X"00000000";
		ram_buffer(15515) := X"00000000";
		ram_buffer(15516) := X"00000000";
		ram_buffer(15517) := X"00000000";
		ram_buffer(15518) := X"00000000";
		ram_buffer(15519) := X"00000000";
		ram_buffer(15520) := X"00000000";
		ram_buffer(15521) := X"00000000";
		ram_buffer(15522) := X"00000000";
		ram_buffer(15523) := X"00000000";
		ram_buffer(15524) := X"00000000";
		ram_buffer(15525) := X"00000000";
		ram_buffer(15526) := X"00000000";
		ram_buffer(15527) := X"00000000";
		ram_buffer(15528) := X"00000000";
		ram_buffer(15529) := X"00000000";
		ram_buffer(15530) := X"00000000";
		ram_buffer(15531) := X"00000000";
		ram_buffer(15532) := X"00000000";
		ram_buffer(15533) := X"00000000";
		ram_buffer(15534) := X"00000000";
		ram_buffer(15535) := X"00000000";
		ram_buffer(15536) := X"00000000";
		ram_buffer(15537) := X"00000000";
		ram_buffer(15538) := X"00000000";
		ram_buffer(15539) := X"00000000";
		ram_buffer(15540) := X"00000000";
		ram_buffer(15541) := X"00000000";
		ram_buffer(15542) := X"00000000";
		ram_buffer(15543) := X"00000000";
		ram_buffer(15544) := X"00000000";
		ram_buffer(15545) := X"00000000";
		ram_buffer(15546) := X"00000000";
		ram_buffer(15547) := X"00000000";
		ram_buffer(15548) := X"00000000";
		ram_buffer(15549) := X"00000000";
		ram_buffer(15550) := X"00000000";
		ram_buffer(15551) := X"00000000";
		ram_buffer(15552) := X"00000000";
		ram_buffer(15553) := X"00000000";
		ram_buffer(15554) := X"00000000";
		ram_buffer(15555) := X"00000000";
		ram_buffer(15556) := X"00000000";
		ram_buffer(15557) := X"00000000";
		ram_buffer(15558) := X"00000000";
		ram_buffer(15559) := X"00000000";
		ram_buffer(15560) := X"00000000";
		ram_buffer(15561) := X"00000000";
		ram_buffer(15562) := X"00000000";
		ram_buffer(15563) := X"00000000";
		ram_buffer(15564) := X"00000000";
		ram_buffer(15565) := X"00000000";
		ram_buffer(15566) := X"00000000";
		ram_buffer(15567) := X"00000000";
		ram_buffer(15568) := X"00000000";
		ram_buffer(15569) := X"00000000";
		ram_buffer(15570) := X"00000000";
		ram_buffer(15571) := X"00000000";
		ram_buffer(15572) := X"00000000";
		ram_buffer(15573) := X"00000000";
		ram_buffer(15574) := X"00000000";
		ram_buffer(15575) := X"00000000";
		ram_buffer(15576) := X"00000000";
		ram_buffer(15577) := X"00000000";
		ram_buffer(15578) := X"00000000";
		ram_buffer(15579) := X"00000000";
		ram_buffer(15580) := X"00000000";
		ram_buffer(15581) := X"00000000";
		ram_buffer(15582) := X"00000000";
		ram_buffer(15583) := X"00000000";
		ram_buffer(15584) := X"00000000";
		ram_buffer(15585) := X"00000000";
		ram_buffer(15586) := X"00000000";
		ram_buffer(15587) := X"00000000";
		ram_buffer(15588) := X"00000000";
		ram_buffer(15589) := X"00000000";
		ram_buffer(15590) := X"00000000";
		ram_buffer(15591) := X"00000000";
		ram_buffer(15592) := X"00000000";
		ram_buffer(15593) := X"00000000";
		ram_buffer(15594) := X"00000000";
		ram_buffer(15595) := X"00000000";
		ram_buffer(15596) := X"00000000";
		ram_buffer(15597) := X"00000000";
		ram_buffer(15598) := X"00000000";
		ram_buffer(15599) := X"00000000";
		ram_buffer(15600) := X"00000000";
		ram_buffer(15601) := X"00000000";
		ram_buffer(15602) := X"00000000";
		ram_buffer(15603) := X"00000000";
		ram_buffer(15604) := X"00000000";
		ram_buffer(15605) := X"00000000";
		ram_buffer(15606) := X"00000000";
		ram_buffer(15607) := X"00000000";
		ram_buffer(15608) := X"00000000";
		ram_buffer(15609) := X"00000000";
		ram_buffer(15610) := X"00000000";
		ram_buffer(15611) := X"00000000";
		ram_buffer(15612) := X"00000000";
		ram_buffer(15613) := X"00000000";
		ram_buffer(15614) := X"00000000";
		ram_buffer(15615) := X"00000000";
		ram_buffer(15616) := X"00000000";
		ram_buffer(15617) := X"00000000";
		ram_buffer(15618) := X"00000000";
		ram_buffer(15619) := X"00000000";
		ram_buffer(15620) := X"00000000";
		ram_buffer(15621) := X"00000000";
		ram_buffer(15622) := X"00000000";
		ram_buffer(15623) := X"00000000";
		ram_buffer(15624) := X"00000000";
		ram_buffer(15625) := X"00000000";
		ram_buffer(15626) := X"00000000";
		ram_buffer(15627) := X"00000000";
		ram_buffer(15628) := X"00000000";
		ram_buffer(15629) := X"00000000";
		ram_buffer(15630) := X"00000000";
		ram_buffer(15631) := X"00000000";
		ram_buffer(15632) := X"00000000";
		ram_buffer(15633) := X"00000000";
		ram_buffer(15634) := X"00000000";
		ram_buffer(15635) := X"00000000";
		ram_buffer(15636) := X"00000000";
		ram_buffer(15637) := X"00000000";
		ram_buffer(15638) := X"00000000";
		ram_buffer(15639) := X"00000000";
		ram_buffer(15640) := X"00000000";
		ram_buffer(15641) := X"00000000";
		ram_buffer(15642) := X"00000000";
		ram_buffer(15643) := X"00000000";
		ram_buffer(15644) := X"00000000";
		ram_buffer(15645) := X"00000000";
		ram_buffer(15646) := X"00000000";
		ram_buffer(15647) := X"00000000";
		ram_buffer(15648) := X"00000000";
		ram_buffer(15649) := X"00000000";
		ram_buffer(15650) := X"00000000";
		ram_buffer(15651) := X"00000000";
		ram_buffer(15652) := X"00000000";
		ram_buffer(15653) := X"00000000";
		ram_buffer(15654) := X"00000000";
		ram_buffer(15655) := X"00000000";
		ram_buffer(15656) := X"00000000";
		ram_buffer(15657) := X"00000000";
		ram_buffer(15658) := X"00000000";
		ram_buffer(15659) := X"00000000";
		ram_buffer(15660) := X"00000000";
		ram_buffer(15661) := X"00000000";
		ram_buffer(15662) := X"00000000";
		ram_buffer(15663) := X"00000000";
		ram_buffer(15664) := X"00000000";
		ram_buffer(15665) := X"00000000";
		ram_buffer(15666) := X"00000000";
		ram_buffer(15667) := X"00000000";
		ram_buffer(15668) := X"00000000";
		ram_buffer(15669) := X"00000000";
		ram_buffer(15670) := X"00000000";
		ram_buffer(15671) := X"00000000";
		ram_buffer(15672) := X"00000000";
		ram_buffer(15673) := X"00000000";
		ram_buffer(15674) := X"00000000";
		ram_buffer(15675) := X"00000000";
		ram_buffer(15676) := X"00000000";
		ram_buffer(15677) := X"00000000";
		ram_buffer(15678) := X"00000000";
		ram_buffer(15679) := X"00000000";
		ram_buffer(15680) := X"00000000";
		ram_buffer(15681) := X"00000000";
		ram_buffer(15682) := X"00000000";
		ram_buffer(15683) := X"00000000";
		ram_buffer(15684) := X"00000000";
		ram_buffer(15685) := X"00000000";
		ram_buffer(15686) := X"00000000";
		ram_buffer(15687) := X"00000000";
		ram_buffer(15688) := X"00000000";
		ram_buffer(15689) := X"00000000";
		ram_buffer(15690) := X"00000000";
		ram_buffer(15691) := X"00000000";
		ram_buffer(15692) := X"00000000";
		ram_buffer(15693) := X"00000000";
		ram_buffer(15694) := X"00000000";
		ram_buffer(15695) := X"00000000";
		ram_buffer(15696) := X"00000000";
		ram_buffer(15697) := X"00000000";
		ram_buffer(15698) := X"00000000";
		ram_buffer(15699) := X"00000000";
		ram_buffer(15700) := X"00000000";
		ram_buffer(15701) := X"00000000";
		ram_buffer(15702) := X"00000000";
		ram_buffer(15703) := X"00000000";
		ram_buffer(15704) := X"00000000";
		ram_buffer(15705) := X"00000000";
		ram_buffer(15706) := X"00000000";
		ram_buffer(15707) := X"00000000";
		ram_buffer(15708) := X"00000000";
		ram_buffer(15709) := X"00000000";
		ram_buffer(15710) := X"00000000";
		ram_buffer(15711) := X"00000000";
		ram_buffer(15712) := X"00000000";
		ram_buffer(15713) := X"00000000";
		ram_buffer(15714) := X"00000000";
		ram_buffer(15715) := X"00000000";
		ram_buffer(15716) := X"00000000";
		ram_buffer(15717) := X"00000000";
		ram_buffer(15718) := X"00000000";
		ram_buffer(15719) := X"00000000";
		ram_buffer(15720) := X"00000000";
		ram_buffer(15721) := X"00000000";
		ram_buffer(15722) := X"00000000";
		ram_buffer(15723) := X"00000000";
		ram_buffer(15724) := X"00000000";
		ram_buffer(15725) := X"00000000";
		ram_buffer(15726) := X"00000000";
		ram_buffer(15727) := X"00000000";
		ram_buffer(15728) := X"00000000";
		ram_buffer(15729) := X"00000000";
		ram_buffer(15730) := X"00000000";
		ram_buffer(15731) := X"00000000";
		ram_buffer(15732) := X"00000000";
		ram_buffer(15733) := X"00000000";
		ram_buffer(15734) := X"00000000";
		ram_buffer(15735) := X"00000000";
		ram_buffer(15736) := X"00000000";
		ram_buffer(15737) := X"00000000";
		ram_buffer(15738) := X"00000000";
		ram_buffer(15739) := X"00000000";
		ram_buffer(15740) := X"00000000";
		ram_buffer(15741) := X"00000000";
		ram_buffer(15742) := X"00000000";
		ram_buffer(15743) := X"00000000";
		ram_buffer(15744) := X"00000000";
		ram_buffer(15745) := X"00000000";
		ram_buffer(15746) := X"00000000";
		ram_buffer(15747) := X"00000000";
		ram_buffer(15748) := X"00000000";
		ram_buffer(15749) := X"00000000";
		ram_buffer(15750) := X"00000000";
		ram_buffer(15751) := X"00000000";
		ram_buffer(15752) := X"00000000";
		ram_buffer(15753) := X"00000000";
		ram_buffer(15754) := X"00000000";
		ram_buffer(15755) := X"00000000";
		ram_buffer(15756) := X"00000000";
		ram_buffer(15757) := X"00000000";
		ram_buffer(15758) := X"00000000";
		ram_buffer(15759) := X"00000000";
		ram_buffer(15760) := X"00000000";
		ram_buffer(15761) := X"00000000";
		ram_buffer(15762) := X"00000000";
		ram_buffer(15763) := X"00000000";
		ram_buffer(15764) := X"00000000";
		ram_buffer(15765) := X"00000000";
		ram_buffer(15766) := X"00000000";
		ram_buffer(15767) := X"00000000";
		ram_buffer(15768) := X"00000000";
		ram_buffer(15769) := X"00000000";
		ram_buffer(15770) := X"00000000";
		ram_buffer(15771) := X"00000000";
		ram_buffer(15772) := X"00000000";
		ram_buffer(15773) := X"00000000";
		ram_buffer(15774) := X"00000000";
		ram_buffer(15775) := X"00000000";
		ram_buffer(15776) := X"00000000";
		ram_buffer(15777) := X"00000000";
		ram_buffer(15778) := X"00000000";
		ram_buffer(15779) := X"00000000";
		ram_buffer(15780) := X"00000000";
		ram_buffer(15781) := X"00000000";
		ram_buffer(15782) := X"00000000";
		ram_buffer(15783) := X"00000000";
		ram_buffer(15784) := X"00000000";
		ram_buffer(15785) := X"00000000";
		ram_buffer(15786) := X"00000000";
		ram_buffer(15787) := X"00000000";
		ram_buffer(15788) := X"00000000";
		ram_buffer(15789) := X"00000000";
		ram_buffer(15790) := X"00000000";
		ram_buffer(15791) := X"00000000";
		ram_buffer(15792) := X"00000000";
		ram_buffer(15793) := X"00000000";
		ram_buffer(15794) := X"00000000";
		ram_buffer(15795) := X"00000000";
		ram_buffer(15796) := X"00000000";
		ram_buffer(15797) := X"00000000";
		ram_buffer(15798) := X"00000000";
		ram_buffer(15799) := X"00000000";
		ram_buffer(15800) := X"00000000";
		ram_buffer(15801) := X"00000000";
		ram_buffer(15802) := X"00000000";
		ram_buffer(15803) := X"00000000";
		ram_buffer(15804) := X"00000000";
		ram_buffer(15805) := X"00000000";
		ram_buffer(15806) := X"00000000";
		ram_buffer(15807) := X"00000000";
		ram_buffer(15808) := X"00000000";
		ram_buffer(15809) := X"00000000";
		ram_buffer(15810) := X"00000000";
		ram_buffer(15811) := X"00000000";
		ram_buffer(15812) := X"00000000";
		ram_buffer(15813) := X"00000000";
		ram_buffer(15814) := X"00000000";
		ram_buffer(15815) := X"00000000";
		ram_buffer(15816) := X"00000000";
		ram_buffer(15817) := X"00000000";
		ram_buffer(15818) := X"00000000";
		ram_buffer(15819) := X"00000000";
		ram_buffer(15820) := X"00000000";
		ram_buffer(15821) := X"00000000";
		ram_buffer(15822) := X"00000000";
		ram_buffer(15823) := X"00000000";
		ram_buffer(15824) := X"00000000";
		ram_buffer(15825) := X"00000000";
		ram_buffer(15826) := X"00000000";
		ram_buffer(15827) := X"00000000";
		ram_buffer(15828) := X"00000000";
		ram_buffer(15829) := X"00000000";
		ram_buffer(15830) := X"00000000";
		ram_buffer(15831) := X"00000000";
		ram_buffer(15832) := X"00000000";
		ram_buffer(15833) := X"00000000";
		ram_buffer(15834) := X"00000000";
		ram_buffer(15835) := X"00000000";
		ram_buffer(15836) := X"00000000";
		ram_buffer(15837) := X"00000000";
		ram_buffer(15838) := X"00000000";
		ram_buffer(15839) := X"00000000";
		ram_buffer(15840) := X"00000000";
		ram_buffer(15841) := X"00000000";
		ram_buffer(15842) := X"00000000";
		ram_buffer(15843) := X"00000000";
		ram_buffer(15844) := X"00000000";
		ram_buffer(15845) := X"00000000";
		ram_buffer(15846) := X"00000000";
		ram_buffer(15847) := X"00000000";
		ram_buffer(15848) := X"00000000";
		ram_buffer(15849) := X"00000000";
		ram_buffer(15850) := X"00000000";
		ram_buffer(15851) := X"00000000";
		ram_buffer(15852) := X"00000000";
		ram_buffer(15853) := X"00000000";
		ram_buffer(15854) := X"00000000";
		ram_buffer(15855) := X"00000000";
		ram_buffer(15856) := X"00000000";
		ram_buffer(15857) := X"00000000";
		ram_buffer(15858) := X"00000000";
		ram_buffer(15859) := X"00000000";
		ram_buffer(15860) := X"00000000";
		ram_buffer(15861) := X"00000000";
		ram_buffer(15862) := X"00000000";
		ram_buffer(15863) := X"00000000";
		ram_buffer(15864) := X"00000000";
		ram_buffer(15865) := X"00000000";
		ram_buffer(15866) := X"00000000";
		ram_buffer(15867) := X"00000000";
		ram_buffer(15868) := X"00000000";
		ram_buffer(15869) := X"00000000";
		ram_buffer(15870) := X"00000000";
		ram_buffer(15871) := X"00000000";
		ram_buffer(15872) := X"00000000";
		ram_buffer(15873) := X"00000000";
		ram_buffer(15874) := X"00000000";
		ram_buffer(15875) := X"00000000";
		ram_buffer(15876) := X"00000000";
		ram_buffer(15877) := X"00000000";
		ram_buffer(15878) := X"00000000";
		ram_buffer(15879) := X"00000000";
		ram_buffer(15880) := X"00000000";
		ram_buffer(15881) := X"00000000";
		ram_buffer(15882) := X"00000000";
		ram_buffer(15883) := X"00000000";
		ram_buffer(15884) := X"00000000";
		ram_buffer(15885) := X"00000000";
		ram_buffer(15886) := X"00000000";
		ram_buffer(15887) := X"00000000";
		ram_buffer(15888) := X"00000000";
		ram_buffer(15889) := X"00000000";
		ram_buffer(15890) := X"00000000";
		ram_buffer(15891) := X"00000000";
		ram_buffer(15892) := X"00000000";
		ram_buffer(15893) := X"00000000";
		ram_buffer(15894) := X"00000000";
		ram_buffer(15895) := X"00000000";
		ram_buffer(15896) := X"00000000";
		ram_buffer(15897) := X"00000000";
		ram_buffer(15898) := X"00000000";
		ram_buffer(15899) := X"00000000";
		ram_buffer(15900) := X"00000000";
		ram_buffer(15901) := X"00000000";
		ram_buffer(15902) := X"00000000";
		ram_buffer(15903) := X"00000000";
		ram_buffer(15904) := X"00000000";
		ram_buffer(15905) := X"00000000";
		ram_buffer(15906) := X"00000000";
		ram_buffer(15907) := X"00000000";
		ram_buffer(15908) := X"00000000";
		ram_buffer(15909) := X"00000000";
		ram_buffer(15910) := X"00000000";
		ram_buffer(15911) := X"00000000";
		ram_buffer(15912) := X"00000000";
		ram_buffer(15913) := X"00000000";
		ram_buffer(15914) := X"00000000";
		ram_buffer(15915) := X"00000000";
		ram_buffer(15916) := X"00000000";
		ram_buffer(15917) := X"00000000";
		ram_buffer(15918) := X"00000000";
		ram_buffer(15919) := X"00000000";
		ram_buffer(15920) := X"00000000";
		ram_buffer(15921) := X"00000000";
		ram_buffer(15922) := X"00000000";
		ram_buffer(15923) := X"00000000";
		ram_buffer(15924) := X"00000000";
		ram_buffer(15925) := X"00000000";
		ram_buffer(15926) := X"00000000";
		ram_buffer(15927) := X"00000000";
		ram_buffer(15928) := X"00000000";
		ram_buffer(15929) := X"00000000";
		ram_buffer(15930) := X"00000000";
		ram_buffer(15931) := X"00000000";
		ram_buffer(15932) := X"00000000";
		ram_buffer(15933) := X"00000000";
		ram_buffer(15934) := X"00000000";
		ram_buffer(15935) := X"00000000";
		ram_buffer(15936) := X"00000000";
		ram_buffer(15937) := X"00000000";
		ram_buffer(15938) := X"00000000";
		ram_buffer(15939) := X"00000000";
		ram_buffer(15940) := X"00000000";
		ram_buffer(15941) := X"00000000";
		ram_buffer(15942) := X"00000000";
		ram_buffer(15943) := X"00000000";
		ram_buffer(15944) := X"00000000";
		ram_buffer(15945) := X"00000000";
		ram_buffer(15946) := X"00000000";
		ram_buffer(15947) := X"00000000";
		ram_buffer(15948) := X"00000000";
		ram_buffer(15949) := X"00000000";
		ram_buffer(15950) := X"00000000";
		ram_buffer(15951) := X"00000000";
		ram_buffer(15952) := X"00000000";
		ram_buffer(15953) := X"00000000";
		ram_buffer(15954) := X"00000000";
		ram_buffer(15955) := X"00000000";
		ram_buffer(15956) := X"00000000";
		ram_buffer(15957) := X"00000000";
		ram_buffer(15958) := X"00000000";
		ram_buffer(15959) := X"00000000";
		ram_buffer(15960) := X"00000000";
		ram_buffer(15961) := X"00000000";
		ram_buffer(15962) := X"00000000";
		ram_buffer(15963) := X"00000000";
		ram_buffer(15964) := X"00000000";
		ram_buffer(15965) := X"00000000";
		ram_buffer(15966) := X"00000000";
		ram_buffer(15967) := X"00000000";
		ram_buffer(15968) := X"00000000";
		ram_buffer(15969) := X"00000000";
		ram_buffer(15970) := X"00000000";
		ram_buffer(15971) := X"00000000";
		ram_buffer(15972) := X"00000000";
		ram_buffer(15973) := X"00000000";
		ram_buffer(15974) := X"00000000";
		ram_buffer(15975) := X"00000000";
		ram_buffer(15976) := X"00000000";
		ram_buffer(15977) := X"00000000";
		ram_buffer(15978) := X"00000000";
		ram_buffer(15979) := X"00000000";
		ram_buffer(15980) := X"00000000";
		ram_buffer(15981) := X"00000000";
		ram_buffer(15982) := X"00000000";
		ram_buffer(15983) := X"00000000";
		ram_buffer(15984) := X"00000000";
		ram_buffer(15985) := X"00000000";
		ram_buffer(15986) := X"00000000";
		ram_buffer(15987) := X"00000000";
		ram_buffer(15988) := X"00000000";
		ram_buffer(15989) := X"00000000";
		ram_buffer(15990) := X"00000000";
		ram_buffer(15991) := X"00000000";
		ram_buffer(15992) := X"00000000";
		ram_buffer(15993) := X"00000000";
		ram_buffer(15994) := X"00000000";
		ram_buffer(15995) := X"00000000";
		ram_buffer(15996) := X"00000000";
		ram_buffer(15997) := X"00000000";
		ram_buffer(15998) := X"00000000";
		ram_buffer(15999) := X"00000000";
		ram_buffer(16000) := X"00000000";
		ram_buffer(16001) := X"00000000";
		ram_buffer(16002) := X"00000000";
		ram_buffer(16003) := X"00000000";
		ram_buffer(16004) := X"00000000";
		ram_buffer(16005) := X"00000000";
		ram_buffer(16006) := X"00000000";
		ram_buffer(16007) := X"00000000";
		ram_buffer(16008) := X"00000000";
		ram_buffer(16009) := X"00000000";
		ram_buffer(16010) := X"00000000";
		ram_buffer(16011) := X"00000000";
		ram_buffer(16012) := X"00000000";
		ram_buffer(16013) := X"00000000";
		ram_buffer(16014) := X"00000000";
		ram_buffer(16015) := X"00000000";
		ram_buffer(16016) := X"00000000";
		ram_buffer(16017) := X"00000000";
		ram_buffer(16018) := X"00000000";
		ram_buffer(16019) := X"00000000";
		ram_buffer(16020) := X"00000000";
		ram_buffer(16021) := X"00000000";
		ram_buffer(16022) := X"00000000";
		ram_buffer(16023) := X"00000000";
		ram_buffer(16024) := X"00000000";
		ram_buffer(16025) := X"00000000";
		ram_buffer(16026) := X"00000000";
		ram_buffer(16027) := X"00000000";
		ram_buffer(16028) := X"00000000";
		ram_buffer(16029) := X"00000000";
		ram_buffer(16030) := X"00000000";
		ram_buffer(16031) := X"00000000";
		ram_buffer(16032) := X"00000000";
		ram_buffer(16033) := X"00000000";
		ram_buffer(16034) := X"00000000";
		ram_buffer(16035) := X"00000000";
		ram_buffer(16036) := X"00000000";
		ram_buffer(16037) := X"00000000";
		ram_buffer(16038) := X"00000000";
		ram_buffer(16039) := X"00000000";
		ram_buffer(16040) := X"00000000";
		ram_buffer(16041) := X"00000000";
		ram_buffer(16042) := X"00000000";
		ram_buffer(16043) := X"00000000";
		ram_buffer(16044) := X"00000000";
		ram_buffer(16045) := X"00000000";
		ram_buffer(16046) := X"00000000";
		ram_buffer(16047) := X"00000000";
		ram_buffer(16048) := X"00000000";
		ram_buffer(16049) := X"00000000";
		ram_buffer(16050) := X"00000000";
		ram_buffer(16051) := X"00000000";
		ram_buffer(16052) := X"00000000";
		ram_buffer(16053) := X"00000000";
		ram_buffer(16054) := X"00000000";
		ram_buffer(16055) := X"00000000";
		ram_buffer(16056) := X"00000000";
		ram_buffer(16057) := X"00000000";
		ram_buffer(16058) := X"00000000";
		ram_buffer(16059) := X"00000000";
		ram_buffer(16060) := X"00000000";
		ram_buffer(16061) := X"00000000";
		ram_buffer(16062) := X"00000000";
		ram_buffer(16063) := X"00000000";
		ram_buffer(16064) := X"00000000";
		ram_buffer(16065) := X"00000000";
		ram_buffer(16066) := X"00000000";
		ram_buffer(16067) := X"00000000";
		ram_buffer(16068) := X"00000000";
		ram_buffer(16069) := X"00000000";
		ram_buffer(16070) := X"00000000";
		ram_buffer(16071) := X"00000000";
		ram_buffer(16072) := X"00000000";
		ram_buffer(16073) := X"00000000";
		ram_buffer(16074) := X"00000000";
		ram_buffer(16075) := X"00000000";
		ram_buffer(16076) := X"00000000";
		ram_buffer(16077) := X"00000000";
		ram_buffer(16078) := X"00000000";
		ram_buffer(16079) := X"00000000";
		ram_buffer(16080) := X"00000000";
		ram_buffer(16081) := X"00000000";
		ram_buffer(16082) := X"00000000";
		ram_buffer(16083) := X"00000000";
		ram_buffer(16084) := X"00000000";
		ram_buffer(16085) := X"00000000";
		ram_buffer(16086) := X"00000000";
		ram_buffer(16087) := X"00000000";
		ram_buffer(16088) := X"00000000";
		ram_buffer(16089) := X"00000000";
		ram_buffer(16090) := X"00000000";
		ram_buffer(16091) := X"00000000";
		ram_buffer(16092) := X"00000000";
		ram_buffer(16093) := X"00000000";
		ram_buffer(16094) := X"00000000";
		ram_buffer(16095) := X"00000000";
		ram_buffer(16096) := X"00000000";
		ram_buffer(16097) := X"00000000";
		ram_buffer(16098) := X"00000000";
		ram_buffer(16099) := X"00000000";
		ram_buffer(16100) := X"00000000";
		ram_buffer(16101) := X"00000000";
		ram_buffer(16102) := X"00000000";
		ram_buffer(16103) := X"00000000";
		ram_buffer(16104) := X"00000000";
		ram_buffer(16105) := X"00000000";
		ram_buffer(16106) := X"00000000";
		ram_buffer(16107) := X"00000000";
		ram_buffer(16108) := X"00000000";
		ram_buffer(16109) := X"00000000";
		ram_buffer(16110) := X"00000000";
		ram_buffer(16111) := X"00000000";
		ram_buffer(16112) := X"00000000";
		ram_buffer(16113) := X"00000000";
		ram_buffer(16114) := X"00000000";
		ram_buffer(16115) := X"00000000";
		ram_buffer(16116) := X"00000000";
		ram_buffer(16117) := X"00000000";
		ram_buffer(16118) := X"00000000";
		ram_buffer(16119) := X"00000000";
		ram_buffer(16120) := X"00000000";
		ram_buffer(16121) := X"00000000";
		ram_buffer(16122) := X"00000000";
		ram_buffer(16123) := X"00000000";
		ram_buffer(16124) := X"00000000";
		ram_buffer(16125) := X"00000000";
		ram_buffer(16126) := X"00000000";
		ram_buffer(16127) := X"00000000";
		ram_buffer(16128) := X"00000000";
		ram_buffer(16129) := X"00000000";
		ram_buffer(16130) := X"00000000";
		ram_buffer(16131) := X"00000000";
		ram_buffer(16132) := X"00000000";
		ram_buffer(16133) := X"00000000";
		ram_buffer(16134) := X"00000000";
		ram_buffer(16135) := X"00000000";
		ram_buffer(16136) := X"00000000";
		ram_buffer(16137) := X"00000000";
		ram_buffer(16138) := X"00000000";
		ram_buffer(16139) := X"00000000";
		ram_buffer(16140) := X"00000000";
		ram_buffer(16141) := X"00000000";
		ram_buffer(16142) := X"00000000";
		ram_buffer(16143) := X"00000000";
		ram_buffer(16144) := X"00000000";
		ram_buffer(16145) := X"00000000";
		ram_buffer(16146) := X"00000000";
		ram_buffer(16147) := X"00000000";
		ram_buffer(16148) := X"00000000";
		ram_buffer(16149) := X"00000000";
		ram_buffer(16150) := X"00000000";
		ram_buffer(16151) := X"00000000";
		ram_buffer(16152) := X"00000000";
		ram_buffer(16153) := X"00000000";
		ram_buffer(16154) := X"00000000";
		ram_buffer(16155) := X"00000000";
		ram_buffer(16156) := X"00000000";
		ram_buffer(16157) := X"00000000";
		ram_buffer(16158) := X"00000000";
		ram_buffer(16159) := X"00000000";
		ram_buffer(16160) := X"00000000";
		ram_buffer(16161) := X"00000000";
		ram_buffer(16162) := X"00000000";
		ram_buffer(16163) := X"00000000";
		ram_buffer(16164) := X"00000000";
		ram_buffer(16165) := X"00000000";
		ram_buffer(16166) := X"00000000";
		ram_buffer(16167) := X"00000000";
		ram_buffer(16168) := X"00000000";
		ram_buffer(16169) := X"00000000";
		ram_buffer(16170) := X"00000000";
		ram_buffer(16171) := X"00000000";
		ram_buffer(16172) := X"00000000";
		ram_buffer(16173) := X"00000000";
		ram_buffer(16174) := X"00000000";
		ram_buffer(16175) := X"00000000";
		ram_buffer(16176) := X"00000000";
		ram_buffer(16177) := X"00000000";
		ram_buffer(16178) := X"00000000";
		ram_buffer(16179) := X"00000000";
		ram_buffer(16180) := X"00000000";
		ram_buffer(16181) := X"00000000";
		ram_buffer(16182) := X"00000000";
		ram_buffer(16183) := X"00000000";
		ram_buffer(16184) := X"00000000";
		ram_buffer(16185) := X"00000000";
		ram_buffer(16186) := X"00000000";
		ram_buffer(16187) := X"00000000";
		ram_buffer(16188) := X"00000000";
		ram_buffer(16189) := X"00000000";
		ram_buffer(16190) := X"00000000";
		ram_buffer(16191) := X"00000000";
		ram_buffer(16192) := X"00000000";
		ram_buffer(16193) := X"00000000";
		ram_buffer(16194) := X"00000000";
		ram_buffer(16195) := X"00000000";
		ram_buffer(16196) := X"00000000";
		ram_buffer(16197) := X"00000000";
		ram_buffer(16198) := X"00000000";
		ram_buffer(16199) := X"00000000";
		ram_buffer(16200) := X"00000000";
		ram_buffer(16201) := X"00000000";
		ram_buffer(16202) := X"00000000";
		ram_buffer(16203) := X"00000000";
		ram_buffer(16204) := X"00000000";
		ram_buffer(16205) := X"00000000";
		ram_buffer(16206) := X"00000000";
		ram_buffer(16207) := X"00000000";
		ram_buffer(16208) := X"00000000";
		ram_buffer(16209) := X"00000000";
		ram_buffer(16210) := X"00000000";
		ram_buffer(16211) := X"00000000";
		ram_buffer(16212) := X"00000000";
		ram_buffer(16213) := X"00000000";
		ram_buffer(16214) := X"00000000";
		ram_buffer(16215) := X"00000000";
		ram_buffer(16216) := X"00000000";
		ram_buffer(16217) := X"00000000";
		ram_buffer(16218) := X"00000000";
		ram_buffer(16219) := X"00000000";
		ram_buffer(16220) := X"00000000";
		ram_buffer(16221) := X"00000000";
		ram_buffer(16222) := X"00000000";
		ram_buffer(16223) := X"00000000";
		ram_buffer(16224) := X"00000000";
		ram_buffer(16225) := X"00000000";
		ram_buffer(16226) := X"00000000";
		ram_buffer(16227) := X"00000000";
		ram_buffer(16228) := X"00000000";
		ram_buffer(16229) := X"00000000";
		ram_buffer(16230) := X"00000000";
		ram_buffer(16231) := X"00000000";
		ram_buffer(16232) := X"00000000";
		ram_buffer(16233) := X"00000000";
		ram_buffer(16234) := X"00000000";
		ram_buffer(16235) := X"00000000";
		ram_buffer(16236) := X"00000000";
		ram_buffer(16237) := X"00000000";
		ram_buffer(16238) := X"00000000";
		ram_buffer(16239) := X"00000000";
		ram_buffer(16240) := X"00000000";
		ram_buffer(16241) := X"00000000";
		ram_buffer(16242) := X"00000000";
		ram_buffer(16243) := X"00000000";
		ram_buffer(16244) := X"00000000";
		ram_buffer(16245) := X"00000000";
		ram_buffer(16246) := X"00000000";
		ram_buffer(16247) := X"00000000";
		ram_buffer(16248) := X"00000000";
		ram_buffer(16249) := X"00000000";
		ram_buffer(16250) := X"00000000";
		ram_buffer(16251) := X"00000000";
		ram_buffer(16252) := X"00000000";
		ram_buffer(16253) := X"00000000";
		ram_buffer(16254) := X"00000000";
		ram_buffer(16255) := X"00000000";
		ram_buffer(16256) := X"00000000";
		ram_buffer(16257) := X"00000000";
		ram_buffer(16258) := X"00000000";
		ram_buffer(16259) := X"00000000";
		ram_buffer(16260) := X"00000000";
		ram_buffer(16261) := X"00000000";
		ram_buffer(16262) := X"00000000";
		ram_buffer(16263) := X"00000000";
		ram_buffer(16264) := X"00000000";
		ram_buffer(16265) := X"00000000";
		ram_buffer(16266) := X"00000000";
		ram_buffer(16267) := X"00000000";
		ram_buffer(16268) := X"00000000";
		ram_buffer(16269) := X"00000000";
		ram_buffer(16270) := X"00000000";
		ram_buffer(16271) := X"00000000";
		ram_buffer(16272) := X"00000000";
		ram_buffer(16273) := X"00000000";
		ram_buffer(16274) := X"00000000";
		ram_buffer(16275) := X"00000000";
		ram_buffer(16276) := X"00000000";
		ram_buffer(16277) := X"00000000";
		ram_buffer(16278) := X"00000000";
		ram_buffer(16279) := X"00000000";
		ram_buffer(16280) := X"00000000";
		ram_buffer(16281) := X"00000000";
		ram_buffer(16282) := X"00000000";
		ram_buffer(16283) := X"00000000";
		ram_buffer(16284) := X"00000000";
		ram_buffer(16285) := X"00000000";
		ram_buffer(16286) := X"00000000";
		ram_buffer(16287) := X"00000000";
		ram_buffer(16288) := X"00000000";
		ram_buffer(16289) := X"00000000";
		ram_buffer(16290) := X"00000000";
		ram_buffer(16291) := X"00000000";
		ram_buffer(16292) := X"00000000";
		ram_buffer(16293) := X"00000000";
		ram_buffer(16294) := X"00000000";
		ram_buffer(16295) := X"00000000";
		ram_buffer(16296) := X"00000000";
		ram_buffer(16297) := X"00000000";
		ram_buffer(16298) := X"00000000";
		ram_buffer(16299) := X"00000000";
		ram_buffer(16300) := X"00000000";
		ram_buffer(16301) := X"00000000";
		ram_buffer(16302) := X"00000000";
		ram_buffer(16303) := X"00000000";
		ram_buffer(16304) := X"00000000";
		ram_buffer(16305) := X"00000000";
		ram_buffer(16306) := X"00000000";
		ram_buffer(16307) := X"00000000";
		ram_buffer(16308) := X"00000000";
		ram_buffer(16309) := X"00000000";
		ram_buffer(16310) := X"00000000";
		ram_buffer(16311) := X"00000000";
		ram_buffer(16312) := X"00000000";
		ram_buffer(16313) := X"00000000";
		ram_buffer(16314) := X"00000000";
		ram_buffer(16315) := X"00000000";
		ram_buffer(16316) := X"00000000";
		ram_buffer(16317) := X"00000000";
		ram_buffer(16318) := X"00000000";
		ram_buffer(16319) := X"00000000";
		ram_buffer(16320) := X"00000000";
		ram_buffer(16321) := X"00000000";
		ram_buffer(16322) := X"00000000";
		ram_buffer(16323) := X"00000000";
		ram_buffer(16324) := X"00000000";
		ram_buffer(16325) := X"00000000";
		ram_buffer(16326) := X"00000000";
		ram_buffer(16327) := X"00000000";
		ram_buffer(16328) := X"00000000";
		ram_buffer(16329) := X"00000000";
		ram_buffer(16330) := X"00000000";
		ram_buffer(16331) := X"00000000";
		ram_buffer(16332) := X"00000000";
		ram_buffer(16333) := X"00000000";
		ram_buffer(16334) := X"00000000";
		ram_buffer(16335) := X"00000000";
		ram_buffer(16336) := X"00000000";
		ram_buffer(16337) := X"00000000";
		ram_buffer(16338) := X"00000000";
		ram_buffer(16339) := X"00000000";
		ram_buffer(16340) := X"00000000";
		ram_buffer(16341) := X"00000000";
		ram_buffer(16342) := X"00000000";
		ram_buffer(16343) := X"00000000";
		ram_buffer(16344) := X"00000000";
		ram_buffer(16345) := X"00000000";
		ram_buffer(16346) := X"00000000";
		ram_buffer(16347) := X"00000000";
		ram_buffer(16348) := X"00000000";
		ram_buffer(16349) := X"00000000";
		ram_buffer(16350) := X"00000000";
		ram_buffer(16351) := X"00000000";
		ram_buffer(16352) := X"00000000";
		ram_buffer(16353) := X"00000000";
		ram_buffer(16354) := X"00000000";
		ram_buffer(16355) := X"00000000";
		ram_buffer(16356) := X"00000000";
		ram_buffer(16357) := X"00000000";
		ram_buffer(16358) := X"00000000";
		ram_buffer(16359) := X"00000000";
		ram_buffer(16360) := X"00000000";
		ram_buffer(16361) := X"00000000";
		ram_buffer(16362) := X"00000000";
		ram_buffer(16363) := X"00000000";
		ram_buffer(16364) := X"00000000";
		ram_buffer(16365) := X"00000000";
		ram_buffer(16366) := X"00000000";
		ram_buffer(16367) := X"00000000";
		ram_buffer(16368) := X"00000000";
		ram_buffer(16369) := X"00000000";
		ram_buffer(16370) := X"00000000";
		ram_buffer(16371) := X"00000000";
		ram_buffer(16372) := X"00000000";
		ram_buffer(16373) := X"00000000";
		ram_buffer(16374) := X"00000000";
		ram_buffer(16375) := X"00000000";
		ram_buffer(16376) := X"00000000";
		ram_buffer(16377) := X"00000000";
		ram_buffer(16378) := X"00000000";
		ram_buffer(16379) := X"00000000";
		ram_buffer(16380) := X"00000000";
		ram_buffer(16381) := X"00000000";
		ram_buffer(16382) := X"00000000";
		ram_buffer(16383) := X"00000000";
		return ram_buffer;
	end;
end;
