memory_initialization_radix=16;
memory_initialization_vector=
3C1C0101,
279CD3B0,
3C050100,
24A553B8,
3C040101,
248457DC,
3C1D0101,
27BD5708,
ACA00000,
00A4182A,
1460FFFD,
24A50004,
0C40007C,
00000000,
0840000E,
23BDFF98,
AFA10010,
AFA20014,
AFA30018,
AFA4001C,
AFA50020,
AFA60024,
AFA70028,
AFA8002C,
AFA90030,
AFAA0034,
AFAB0038,
AFAC003C,
AFAD0040,
AFAE0044,
AFAF0048,
AFB8004C,
AFB90050,
AFBF0054,
401A7000,
235AFFFC,
AFBA0058,
0000D810,
AFBB005C,
0000D812,
AFBB0060,
0C40127B,
23A50000,
8FA10010,
8FA20014,
8FA30018,
8FA4001C,
8FA50020,
8FA60024,
8FA70028,
8FA8002C,
8FA90030,
8FAA0034,
8FAB0038,
8FAC003C,
8FAD0040,
8FAE0044,
8FAF0048,
8FB8004C,
8FB90050,
8FBF0054,
8FBA0058,
8FBB005C,
03600011,
8FBB0060,
03600013,
23BD0068,
341B0001,
03400008,
409B6000,
40026000,
03E00008,
40846000,
3C050100,
24A50150,
8CA60000,
AC06003C,
8CA60004,
AC060040,
8CA60008,
AC060044,
8CA6000C,
03E00008,
AC060048,
3C1A0100,
375A003C,
03400008,
00000000,
AC900000,
AC910004,
AC920008,
AC93000C,
AC940010,
AC950014,
AC960018,
AC97001C,
AC9E0020,
AC9C0024,
AC9D0028,
AC9F002C,
03E00008,
34020000,
8C900000,
8C910004,
8C920008,
8C93000C,
8C940010,
8C950014,
8C960018,
8C97001C,
8C9E0020,
8C9C0024,
8C9D0028,
8C9F002C,
03E00008,
34A20000,
00850019,
00001012,
00002010,
03E00008,
ACC40000,
0000000C,
03E00008,
00000000,
3C040100,
27BDFFE8,
AFBF0014,
0C400256,
248404AC,
8FBF0014,
00001025,
03E00008,
27BD0018,
2082FF78,
AC450078,
03E00008,
AC46001C,
3C1A0100,
375A5420,
8F5B0000,
AF400000,
23BDFF78,
AFA10010,
AFA20014,
AFA30018,
AFA4001C,
AFA50020,
AFA60024,
AFA70028,
AFA8002C,
AFA90030,
AFAA0034,
AFAB0038,
AFAC003C,
AFAD0040,
AFAE0044,
AFAF0048,
AFB0004C,
AFB10050,
AFB20054,
AFB30058,
AFB4005C,
AFB50060,
AFB60064,
AFB70068,
AFB8006C,
AFB90070,
AFBF0074,
401A7000,
17600003,
235AFFFC,
084000AE,
00000000,
235A0004,
AFBA0078,
0000D810,
AFBB007C,
0000D812,
AFBB0080,
3C1A0100,
375A53C8,
8F5A0000,
AF5D0000,
3C1A0101,
375A5520,
8F5D0000,
0C400205,
00000000,
3C1A0101,
375A5520,
AF5D0000,
3C1A0100,
375A53C8,
8F5A0000,
8F5D0000,
8FA10010,
8FA20014,
8FA30018,
8FA4001C,
8FA50020,
8FA60024,
8FA70028,
8FA8002C,
8FA90030,
8FAA0034,
8FAB0038,
8FAC003C,
8FAD0040,
8FAE0044,
8FAF0048,
8FB0004C,
8FB10050,
8FB20054,
8FB30058,
8FB4005C,
8FB50060,
8FB60064,
8FB70068,
8FB8006C,
8FB90070,
8FBF0074,
8FBA0078,
8FBB007C,
03600011,
8FBB0080,
03600013,
23BD0088,
341B0001,
03400008,
409B6000,
00000000,
3C080100,
250803C8,
8D090000,
AC09003C,
8D090004,
AC090040,
8D090008,
AC090044,
8D09000C,
03E00008,
AC090048,
3C1A0100,
375A0224,
03400008,
00000000,
3C1A0101,
375A5520,
AF5D0000,
3C1A0100,
375A53C8,
8F5A0000,
8F5D0000,
8FA10010,
8FA20014,
8FA30018,
8FA4001C,
8FA50020,
8FA60024,
8FA70028,
8FA8002C,
8FA90030,
8FAA0034,
8FAB0038,
8FAC003C,
8FAD0040,
8FAE0044,
8FAF0048,
8FB0004C,
8FB10050,
8FB20054,
8FB30058,
8FB4005C,
8FB50060,
8FB60064,
8FB70068,
8FB8006C,
8FB90070,
8FBF0074,
8FBA0078,
8FBB007C,
03600011,
8FBB0080,
03600013,
23BD0088,
341B0001,
03400008,
409B6000,
40806000,
20090001,
3C080100,
35085420,
AD090000,
3C080100,
35085404,
AD090000,
0000000C,
03E00008,
00000000,
3C060100,
27BDFFE8,
24C60544,
2405001E,
AFBF0014,
0C400288,
00002025,
3C060100,
24C6056C,
24050018,
0C400288,
24040001,
3C060100,
24C6059C,
24050012,
0C400288,
24040002,
3C060100,
24C605CC,
2405000C,
0C400288,
24040003,
3C060100,
24C605FC,
24050006,
0C400288,
24040004,
0C4002A8,
00002025,
3C060100,
24040005,
24C60624,
0C400288,
24050002,
8FBF0014,
24040005,
084002A8,
27BD0018,
27BDFFE8,
AFBF0014,
0C4002A8,
24040001,
8F828084,
00000000,
24420001,
AF828084,
1000FFF9,
00000000,
27BDFFE8,
AFBF0014,
0C4002BE,
24040001,
0C4002A8,
24040002,
8F828080,
00000000,
24420001,
AF828080,
1000FFF7,
00000000,
27BDFFE8,
AFBF0014,
0C4002BE,
24040002,
0C4002A8,
24040003,
8F82807C,
00000000,
24420001,
AF82807C,
1000FFF7,
00000000,
27BDFFE8,
AFBF0014,
0C4002BE,
24040003,
0C4002A8,
24040004,
8F828074,
00000000,
24420001,
AF828074,
1000FFF7,
00000000,
27BDFFE8,
AFBF0014,
0C4002BE,
24040004,
8F828078,
00000000,
24420001,
AF828078,
1000FFF9,
00000000,
27BDFFD0,
AFB40020,
AFB3001C,
AFB10014,
3C130100,
3C140100,
3C110100,
AFB60028,
AFB50024,
AFB20018,
AFBF002C,
AFB00010,
0000A825,
00009025,
26735218,
24160005,
26945260,
263152D0,
2404001E,
0C4002CD,
2652001E,
02402825,
0C4004A5,
02602025,
8F908084,
8F858080,
8F84807C,
02058021,
8F838074,
02048021,
8F828078,
02038021,
02028021,
16C00002,
0216001B,
0007000D,
8F848084,
00001012,
2443FFFF,
0083202B,
1480002E,
00000000,
8F848084,
24420001,
0044202B,
14800029,
00000000,
8F848080,
00000000,
0083202B,
14800024,
00000000,
8F848080,
00000000,
0044202B,
1480001F,
00000000,
8F84807C,
00000000,
0083202B,
1480001A,
00000000,
8F84807C,
00000000,
0044202B,
14800015,
00000000,
8F848074,
00000000,
0083202B,
14800010,
00000000,
8F848074,
00000000,
0044202B,
1480000B,
00000000,
8F848078,
00000000,
0083182B,
14600006,
00000000,
8F838078,
00000000,
0043102B,
10400004,
02152823,
0C4004A5,
02802025,
02152823,
0C4004A5,
02202025,
1000FFB5,
0200A825,
8F838094,
00000000,
8C620000,
00000000,
30420002,
1040FFFC,
00000000,
AC650008,
03E00008,
00000000,
27BDFFE8,
AFBF0014,
0C400A8D,
00000000,
10400002,
24020001,
AF828054,
8FBF0014,
8F82808C,
24030007,
AC430000,
03E00008,
27BD0018,
8F828094,
3C040100,
8C420004,
084004A5,
248452EC,
03E00008,
00000000,
24020001,
3C030101,
AF82800C,
8C625720,
27BDFFE0,
8C420004,
AFB10018,
3C110101,
AFB00014,
AFBF001C,
00608025,
26315724,
2C430008,
14600014,
000210C0,
8F828008,
00000000,
10400004,
00000000,
AF808008,
0C400203,
00000000,
AF80800C,
8F828054,
00000000,
10400012,
00000000,
8FBF001C,
8FB10018,
8FB00014,
27BD0020,
AF808054,
08400B08,
00000000,
02221021,
8C430000,
8C440004,
0060F809,
00000000,
8E025720,
00000000,
8C420004,
1000FFE2,
2C430008,
8FBF001C,
8FB10018,
8FB00014,
03E00008,
27BD0020,
27BDFFE0,
8F828090,
3403FFFF,
AFB00010,
3C100100,
AFB20018,
AFB10014,
AFBF001C,
00808825,
00A09025,
AC430008,
261052F8,
02403025,
02202825,
0C4004A5,
02002025,
1000FFFC,
02403025,
3C020101,
8C425720,
240300FF,
03E00008,
AC430000,
3C020101,
8C425720,
00000000,
03E00008,
AC400000,
24020001,
AF828008,
08400120,
00000000,
27BDFFE8,
AFB00010,
00808025,
AFBF0014,
0C400046,
00002025,
3C0344A0,
3C020101,
AC435720,
3C040101,
3C030101,
24635724,
24845764,
24630008,
1464FFFE,
AC60FFF8,
3C0344A2,
AF838090,
3404C350,
3C0344A1,
AF83808C,
AC640004,
3C030100,
24425720,
246307C4,
AC430004,
3C0344A4,
AF838094,
3C030100,
246307F8,
3C050100,
AC400008,
AC43001C,
AC400020,
24A5079C,
0C4004A2,
00002025,
0200F809,
00000000,
8F82808C,
24030003,
AC430000,
8F828090,
24030001,
0C400D84,
AC430008,
3C040100,
240500CF,
0C400236,
24845318,
00041080,
3C040101,
24845764,
00822021,
2402001F,
00452823,
24020006,
14400002,
00A2001A,
0007000D,
27BDFFE0,
00C01825,
00003825,
AFA40014,
2406012C,
00602025,
AFBF001C,
00002812,
AFA50010,
0C400CC9,
00002825,
24030001,
10430005,
00001025,
3C040100,
240500DD,
0C400236,
24845318,
8FBF001C,
00000000,
03E00008,
27BD0020,
3C030101,
00042080,
24625764,
8F85800C,
27BDFFE8,
00441021,
8C440000,
10A0000A,
AFBF0014,
0C400A24,
00000000,
10400002,
24020001,
AF828054,
8FBF0014,
00001025,
03E00008,
27BD0018,
0C400ED5,
00000000,
1000FFF9,
00000000,
3C020101,
24425764,
00042080,
00822021,
8C840000,
27BDFFE8,
AFBF0014,
0C400E8E,
00000000,
8FBF0014,
00001025,
03E00008,
27BD0018,
08400120,
00000000,
240203E8,
00820018,
00002012,
08400FAD,
00000000,
27BDFFE8,
00003025,
24050010,
AFB00010,
00808025,
24040001,
AFBF0014,
0C4005E6,
00108080,
27848088,
00902021,
14400005,
AC820000,
3C040100,
24050116,
0C400236,
24845318,
8FBF0014,
8FB00010,
00001025,
03E00008,
27BD0018,
8F82800C,
27BDFFE0,
00042080,
10400013,
AFBF001C,
27828088,
00442021,
8C840000,
00003825,
27A60010,
0C400704,
AFA00010,
8FA30010,
00000000,
10600003,
24030001,
AF838054,
24030001,
1043000C,
3C040100,
2405012A,
0C400236,
24845318,
27828088,
00442021,
8C840000,
00003825,
0C400628,
2406FFFF,
1000FFF4,
24030001,
8FBF001C,
00001025,
03E00008,
27BD0020,
8F82800C,
27BDFFE0,
00042080,
10400012,
AFBF001C,
27828088,
00442021,
8C840000,
27A60010,
0C400877,
AFA00010,
8FA30010,
00000000,
10600003,
24030001,
AF838054,
24030001,
1043000C,
3C040100,
2405013E,
0C400236,
24845318,
27828088,
00442021,
8C840000,
00003825,
0C40079E,
2406FFFF,
1000FFF4,
24030001,
8FBF001C,
00001025,
03E00008,
27BD0020,
27BDFFE8,
24050001,
AFB00010,
00808025,
24040001,
AFBF0014,
0C40060A,
00108080,
2784809C,
00902021,
14400005,
AC820000,
3C040100,
2405014A,
0C400236,
24845318,
8FBF0014,
8FB00010,
00001025,
03E00008,
27BD0018,
8F82800C,
27BDFFE0,
00042080,
10400013,
AFBF001C,
2782809C,
00442021,
8C840000,
27A60010,
00002825,
0C400877,
AFA00010,
8FA30010,
00000000,
10600003,
24030001,
AF838054,
24030001,
1043000D,
3C040100,
2405015E,
0C400236,
24845318,
2782809C,
00442021,
8C840000,
00003825,
2406FFFF,
0C40079E,
00002825,
1000FFF3,
24030001,
8FBF001C,
00001025,
03E00008,
27BD0020,
8F82800C,
27BDFFE0,
00042080,
10400012,
AFBF001C,
2782809C,
00442021,
8C840000,
27A50010,
0C40075A,
AFA00010,
8FA30010,
00000000,
10600003,
24030001,
AF838054,
24030001,
1043000D,
3C040100,
24050172,
0C400236,
24845318,
2782809C,
00442021,
8C840000,
00003825,
00003025,
0C400628,
00002825,
1000FFF3,
24030001,
8FBF001C,
00001025,
03E00008,
27BD0020,
03E00008,
00001025,
27BDFFE0,
AFB00014,
00808025,
24040080,
AFB10018,
AFBF001C,
00A08825,
0C4012B1,
00108080,
27848098,
00902021,
AC820000,
14400005,
AE220000,
3C040100,
24050189,
0C400236,
24845318,
8FBF001C,
8FB10018,
8FB00014,
00001025,
03E00008,
27BD0020,
27828098,
00042080,
00442021,
8C840000,
27BDFFE8,
24020001,
14850004,
AFBF0014,
0C401323,
00000000,
00001025,
8FBF0014,
00000000,
03E00008,
27BD0018,
24020001,
14400002,
0082001B,
0007000D,
00001812,
0065182B,
10600006,
00450018,
00004025,
14400006,
00000000,
03E00008,
A0E00000,
00001012,
1000FFF2,
00000000,
14400002,
0082001B,
0007000D,
00002010,
00004812,
00000000,
00000000,
14A00002,
0045001B,
0007000D,
00001012,
15000005,
292A000A,
1D200004,
24EB0001,
1440FFE9,
00000000,
24EB0001,
15400004,
24030030,
14C00002,
24030037,
24030057,
00691821,
A0E30000,
25080001,
1000FFDE,
01603825,
27BDFFD8,
AFB40020,
AFB3001C,
AFB20018,
AFB10014,
AFBF0024,
AFB00010,
00809025,
00A09825,
8FB10038,
10E00002,
24140020,
24140030,
02201025,
24420001,
8043FFFF,
00000000,
14600009,
00C08025,
1A000009,
02802825,
0260F809,
02402025,
1000FFFB,
2610FFFF,
1000FFF4,
24C6FFFF,
1CC0FFFD,
00000000,
26310001,
8225FFFF,
00000000,
14A00009,
00000000,
8FBF0024,
8FB40020,
8FB3001C,
8FB20018,
8FB10014,
8FB00010,
03E00008,
27BD0028,
0260F809,
02402025,
1000FFF1,
26310001,
8C820000,
00000000,
24430001,
AC830000,
03E00008,
A0450000,
27BDFFB8,
AFB5003C,
AFB40038,
AFB30034,
AFB20030,
AFB1002C,
AFB00028,
AFBF0044,
AFB60040,
00809025,
00A09825,
00C08825,
00E08025,
24140025,
24150030,
82250000,
00000000,
10A00035,
00000000,
10B40006,
00000000,
26310001,
0260F809,
02402025,
1000FFF6,
00000000,
82260001,
00000000,
10D50015,
240D0001,
26310002,
00006825,
24C2FFD0,
304200FF,
2C42000A,
10400018,
00006025,
30C200FF,
2443FFD0,
2C63000A,
1060000C,
2443FF9F,
24C3FFD0,
000C1080,
004C6021,
000C6040,
26310001,
8226FFFF,
1000FFF4,
01836021,
82260002,
1000FFEC,
26310003,
2C630006,
1060001A,
2442FFBF,
24C3FFA9,
2862000B,
1440FFF1,
000C1080,
24020063,
10C20045,
28C20064,
10400016,
24020073,
10D4004C,
24020058,
10C20033,
00000000,
14C0FFC9,
00000000,
8FBF0044,
8FB60040,
8FB5003C,
8FB40038,
8FB30034,
8FB20030,
8FB1002C,
8FB00028,
03E00008,
27BD0048,
2C420006,
1040FFEA,
24020063,
1000FFE4,
24C3FFC9,
10C20032,
28C20074,
10400019,
24020075,
24020064,
14C2FFB3,
26160004,
8E040000,
00000000,
04810005,
27A70018,
2402002D,
00042023,
A3A20018,
27A70019,
00003025,
2405000A,
0C4003B2,
00000000,
27A20018,
AFA20010,
01A03825,
01803025,
02602825,
0C4003DE,
02402025,
1000FF9E,
02C08025,
10C2000A,
26160004,
24020078,
14C2FF99,
00000000,
38C60058,
26160004,
27A70018,
2CC60001,
10000004,
24050010,
27A70018,
00003025,
2405000A,
8E040000,
1000FFE5,
00000000,
82050003,
02402025,
0260F809,
26160004,
1000FF87,
02C08025,
8E020000,
26160004,
AFA20010,
1000FFDF,
00003825,
1000FF87,
24050025,
AF858014,
03E00008,
AF848010,
27BDFFE0,
AFA50024,
AFA60028,
8F858014,
00803025,
8F848010,
AFA7002C,
27A70024,
AFBF001C,
0C400412,
AFA70010,
8FBF001C,
00000000,
03E00008,
27BD0020,
27BDFFE0,
AFA60028,
00A03025,
3C050100,
AFA40020,
AFA7002C,
27A40020,
27A70028,
24A51030,
AFBF001C,
0C400412,
AFA70010,
8FA20020,
00000000,
A0400000,
8FBF001C,
00000000,
03E00008,
27BD0020,
10C0000D,
00C53021,
2402FFF0,
00C21824,
0066302B,
00A22824,
00063100,
24620010,
00463021,
3C022000,
00822021,
2402FFF0,
14C50003,
00A21824,
03E00008,
00000000,
AC830000,
AC600000,
1000FFF9,
24A50010,
24820008,
2403FFFF,
AC820004,
AC830008,
AC82000C,
AC820010,
03E00008,
AC800000,
03E00008,
AC800010,
8C820004,
00000000,
8C430008,
ACA20004,
ACA30008,
8C430008,
00000000,
AC650004,
AC450008,
8C820000,
ACA40010,
24420001,
03E00008,
AC820000,
8CA60000,
2403FFFF,
14C3000F,
24820008,
8C820010,
00000000,
8C430004,
00000000,
ACA30004,
AC650008,
ACA20008,
AC450004,
8C820000,
ACA40010,
24420001,
03E00008,
AC820000,
00E01025,
8C470004,
00000000,
8CE30000,
00000000,
00C3182B,
1060FFF9,
00000000,
1000FFEC,
00000000,
8C850004,
8C820008,
8C830010,
ACA20008,
8C820008,
00000000,
AC450004,
8C650004,
00000000,
14850002,
00000000,
AC620004,
8C620000,
AC800010,
2442FFFF,
03E00008,
AC620000,
27BDFFE0,
AFB20018,
00C09025,
8C860040,
AFB10014,
AFB00010,
AFBF001C,
00808025,
8C910038,
14C00011,
00000000,
8C830000,
00000000,
14600005,
00001025,
8C840004,
0C400C61,
00000000,
AE000004,
8FBF001C,
26310001,
AE110038,
8FB20018,
8FB10014,
8FB00010,
03E00008,
27BD0020,
16400010,
00000000,
8C840008,
0C40135C,
00000000,
8E020008,
8E030040,
00000000,
00431021,
8E030004,
AE020008,
0043182B,
1460FFEB,
00001025,
8E030000,
1000FFE8,
AE030008,
8C84000C,
0C40135C,
00000000,
8E030040,
8E02000C,
00031823,
8E040000,
00431021,
AE02000C,
0044102B,
10400005,
00000000,
8E020004,
00000000,
00431821,
AE03000C,
24030002,
1643FFD5,
00001025,
0011182B,
1000FFD2,
02238823,
00801025,
8C460040,
00000000,
10C0000E,
00A02025,
8C43000C,
8C450004,
00661821,
AC43000C,
0065182B,
14600004,
00000000,
8C430000,
00000000,
AC43000C,
8C45000C,
0840135C,
00000000,
03E00008,
00000000,
27BDFFE0,
AFB00010,
AFB20018,
AFB10014,
AFBF001C,
0C400C9C,
00808025,
92110045,
26120024,
00118E00,
00118E03,
1E200013,
2402FFFF,
A2020045,
0C400CAF,
00000000,
0C400C9C,
00000000,
92110044,
26120010,
00118E00,
00118E03,
1E200016,
2402FFFF,
8FBF001C,
8FB20018,
8FB10014,
A2020044,
8FB00010,
08400CAF,
27BD0020,
8E020024,
00000000,
1040FFEB,
2402FFFF,
0C400B7F,
02402025,
10400003,
00000000,
0C400BFF,
00000000,
2631FFFF,
00118E00,
1000FFDF,
00118E03,
8E020010,
00000000,
1040FFE8,
2402FFFF,
0C400B7F,
02402025,
10400003,
00000000,
0C400BFF,
00000000,
2631FFFF,
00118E00,
1000FFDC,
00118E03,
27BDFFE0,
AFB10018,
AFB00014,
AFBF001C,
00808025,
14800005,
00A08825,
3C040100,
2405011B,
0C400236,
24845334,
0C400C9C,
00000000,
8E050040,
8E03003C,
8E040000,
00A30018,
AE000038,
AE040008,
00001012,
00821821,
00451023,
00821021,
AE02000C,
2402FFFF,
A2020044,
AE030004,
A2020045,
16200013,
00000000,
8E020010,
00000000,
10400007,
00000000,
0C400B7F,
26040010,
10400003,
00000000,
0C400120,
00000000,
0C400CAF,
00000000,
8FBF001C,
8FB10018,
8FB00014,
24020001,
03E00008,
27BD0020,
0C4004DB,
26040010,
0C4004DB,
26040024,
1000FFF3,
00000000,
27BDFFE0,
AFB20018,
AFB10014,
AFBF001C,
AFB00010,
00809025,
14800005,
00A08825,
3C040100,
24050188,
0C400236,
24845334,
02510018,
00002012,
0C4012B1,
24840048,
10400009,
00408025,
1620000E,
00000000,
AE020000,
AE12003C,
AE110040,
24050001,
0C4005B0,
02002025,
8FBF001C,
02001025,
8FB20018,
8FB10014,
8FB00010,
03E00008,
27BD0020,
24420048,
1000FFF2,
AE020000,
27BDFFE0,
AFB10018,
AFB00014,
AFBF001C,
00808025,
14800005,
00A08825,
3C040100,
240502BD,
0C400236,
24845334,
0211102B,
10400006,
24060002,
3C040100,
240502BE,
0C400236,
24845334,
24060002,
00002825,
0C4005E6,
02002025,
10400002,
00000000,
AC510038,
8FBF001C,
8FB10018,
8FB00014,
03E00008,
27BD0020,
27BDFFC0,
AFB30028,
AFB10020,
AFB0001C,
AFBF003C,
AFB70038,
AFB60034,
AFB50030,
AFB4002C,
AFB20024,
00808025,
00A09825,
AFA60048,
14800005,
00E08825,
3C040100,
240502D9,
0C400236,
24845334,
16600006,
24020002,
8E020040,
00000000,
14400083,
240502DA,
24020002,
16220005,
24020001,
8E03003C,
00000000,
14620081,
3C040100,
0C400C16,
00000000,
14400009,
0000B025,
8FA20048,
00000000,
10400005,
3C040100,
240502DE,
0C400236,
24845334,
0000B025,
24150002,
2412FFFF,
1000003B,
26140010,
8FA20048,
00000000,
14400005,
00000000,
0C400CAF,
00000000,
1000004D,
00001025,
16C00003,
00000000,
0C400BED,
27A40010,
0C400CAF,
00000000,
0C400A61,
00000000,
0C400C9C,
00000000,
92020044,
00000000,
00021600,
00021603,
14520002,
00000000,
A2000044,
92020045,
00000000,
00021600,
00021603,
14520002,
00000000,
A2000045,
0C400CAF,
00000000,
27A50048,
0C401075,
27A40010,
1440003F,
00000000,
0C400C9C,
00000000,
8E170038,
8E16003C,
0C400CAF,
00000000,
16F60031,
00000000,
8FA50048,
0C400B45,
02802025,
0C400575,
02002025,
0C400F0A,
00000000,
14400003,
24160001,
0C400120,
00000000,
0C400C9C,
00000000,
8E020038,
8E03003C,
00000000,
0043102B,
14400003,
02203025,
1635FFBD,
00000000,
02602825,
0C40051F,
02002025,
8E030024,
00000000,
10600003,
00000000,
0C400B7F,
26040024,
10400003,
00000000,
0C400120,
00000000,
0C400CAF,
00000000,
24020001,
8FBF003C,
8FB70038,
8FB60034,
8FB50030,
8FB4002C,
8FB30028,
8FB20024,
8FB10020,
8FB0001C,
03E00008,
27BD0040,
0C400575,
02002025,
0C400F0A,
24160001,
1000FFD6,
00000000,
0C400575,
02002025,
0C400F0A,
00000000,
1000FFEA,
00001025,
3C040100,
0C400236,
24845334,
1000FF7B,
24020002,
240502DB,
0C400236,
24845334,
1000FF7C,
00000000,
27BDFFE8,
00803025,
00002825,
AFB00010,
AFBF0014,
0C4005E6,
24040001,
10400009,
00408025,
AC400004,
AC400000,
AC40000C,
00003825,
00003025,
00002825,
0C400628,
00402025,
8FBF0014,
02001025,
8FB00010,
03E00008,
27BD0018,
27BDFFE0,
AFB00010,
AFBF001C,
AFB20018,
AFB10014,
14800005,
00808025,
3C040100,
24050241,
0C400236,
24845334,
8E120004,
0C400C13,
00008825,
1642000B,
00000000,
8E02000C,
24110001,
2442FFFF,
14400006,
AE02000C,
00003825,
00003025,
00002825,
0C400628,
02002025,
8FBF001C,
02201025,
8FB20018,
8FB10014,
8FB00010,
03E00008,
27BD0020,
27BDFFD0,
AFB40024,
AFB30020,
AFB2001C,
AFB00014,
AFBF002C,
AFB50028,
AFB10018,
00808025,
00A09825,
00C0A025,
14800005,
00E09025,
3C040100,
2405039F,
0C400236,
24845334,
16600006,
24020002,
8E020040,
00000000,
14400036,
240503A0,
24020002,
16420005,
24020001,
8E03003C,
00000000,
14620034,
240503A1,
8E020038,
8E03003C,
00000000,
0043102B,
14400003,
24030002,
16430018,
00000000,
92110045,
02403025,
0011AE00,
02602825,
0C40051F,
02002025,
0015AE03,
2402FFFF,
16A20017,
00000000,
8E020024,
00000000,
14400003,
00000000,
10000008,
24020001,
0C400B7F,
26040024,
1040FFFB,
00000000,
12800002,
24020001,
AE820000,
8FBF002C,
8FB50028,
8FB40024,
8FB30020,
8FB2001C,
8FB10018,
8FB00014,
03E00008,
27BD0030,
26310001,
00118E00,
00118E03,
A2110045,
1000FFF2,
24020001,
3C040100,
0C400236,
24845334,
1000FFC8,
24020002,
3C040100,
0C400236,
24845334,
1000FFC9,
00000000,
27BDFFE0,
AFB10018,
AFB00014,
AFBF001C,
00808025,
14800005,
00A08825,
3C040100,
2405043C,
0C400236,
24845334,
8E020040,
00000000,
10400004,
24050440,
3C040100,
0C400236,
24845334,
8E020000,
00000000,
14400005,
00000000,
8E020004,
00000000,
14400026,
3C040100,
8E030038,
8E04003C,
00000000,
0064202B,
10800016,
00001025,
92020045,
24630001,
00022600,
AE030038,
00042603,
2403FFFF,
14830013,
24420001,
8E020024,
00000000,
14400003,
00000000,
10000008,
24020001,
0C400B7F,
26040024,
1040FFFB,
00000000,
12200002,
24020001,
AE220000,
8FBF001C,
8FB10018,
8FB00014,
03E00008,
27BD0020,
00021600,
00021603,
A2020045,
1000FFF7,
24020001,
24050445,
0C400236,
24845334,
1000FFD7,
00000000,
27BDFFC8,
AFB5002C,
AFB30024,
AFB00018,
AFBF0034,
AFB60030,
AFB40028,
AFB20020,
AFB1001C,
00808025,
00A09825,
AFA60040,
14800005,
00E0A825,
3C040100,
240504DC,
0C400236,
24845334,
16600005,
00000000,
8E020040,
00000000,
14400096,
3C040100,
0C400C16,
00000000,
14400009,
0000B025,
8FA20040,
00000000,
10400005,
3C040100,
240504E0,
0C400236,
24845334,
0000B025,
2412FFFF,
1000004B,
26140024,
8E020024,
AE12000C,
10400063,
26040024,
1000005B,
00000000,
8FA20040,
00000000,
14400005,
00000000,
0C400CAF,
00000000,
1000005C,
00001025,
16C00003,
00000000,
0C400BED,
27A40010,
0C400CAF,
00000000,
0C400A61,
00000000,
0C400C9C,
00000000,
92020044,
00000000,
00021600,
00021603,
14520002,
00000000,
A2000044,
92020045,
00000000,
00021600,
00021603,
14520002,
00000000,
A2000045,
0C400CAF,
00000000,
27A50040,
0C401075,
27A40010,
1440004D,
00000000,
0C400C9C,
00000000,
8E110038,
0C400CAF,
00000000,
16200040,
00000000,
8E020000,
00000000,
14400008,
00000000,
0C400C9C,
00000000,
8E040004,
0C400C20,
00000000,
0C400CAF,
00000000,
8FA50040,
0C400B45,
02802025,
0C400575,
02002025,
0C400F0A,
00000000,
14400003,
24160001,
0C400120,
00000000,
0C400C9C,
00000000,
8E110038,
00000000,
1220FFB7,
02602825,
8E12000C,
0C400561,
02002025,
16A0FFAC,
2631FFFF,
8E020000,
AE110038,
14400004,
00000000,
0C4010BA,
00000000,
AE020004,
8E020010,
00000000,
10400007,
26040010,
0C400B7F,
00000000,
10400003,
00000000,
0C400120,
00000000,
0C400CAF,
00000000,
24020001,
8FBF0034,
8FB60030,
8FB5002C,
8FB40028,
8FB30024,
8FB20020,
8FB1001C,
8FB00018,
03E00008,
27BD0038,
0C400575,
02002025,
0C400F0A,
24160001,
1000FFD2,
00000000,
0C400575,
02002025,
0C400F0A,
00000000,
0C400C9C,
00000000,
8E110038,
0C400CAF,
00000000,
1620FFC7,
24160001,
1000FFE4,
00001025,
240504DD,
0C400236,
24845334,
1000FF67,
00000000,
27BDFFE0,
AFB10014,
AFB00010,
AFBF001C,
AFB20018,
00808025,
14800005,
00A08825,
3C040100,
24050278,
0C400236,
24845334,
8E120004,
0C400C13,
00000000,
1642000C,
00003825,
8E02000C,
00000000,
24420001,
AE02000C,
24020001,
8FBF001C,
8FB20018,
8FB10014,
8FB00010,
03E00008,
27BD0020,
02203025,
00002825,
0C40079E,
02002025,
1040FFF5,
00000000,
8E03000C,
00000000,
24630001,
1000FFF0,
AE03000C,
27BDFFD0,
AFB40024,
AFB30020,
AFB00014,
AFBF002C,
AFB50028,
AFB2001C,
AFB10018,
00808025,
00A09825,
14800005,
00C0A025,
3C040100,
240505A0,
0C400236,
24845334,
16600005,
00000000,
8E020040,
00000000,
1440002C,
240505A1,
8E120038,
00000000,
12400019,
00001025,
92110044,
02602825,
0011AE00,
0C400561,
02002025,
2652FFFF,
0015AE03,
2402FFFF,
AE120038,
16A20017,
00000000,
8E020010,
00000000,
14400003,
00000000,
10000008,
24020001,
0C400B7F,
26040010,
1040FFFB,
00000000,
12800002,
24020001,
AE820000,
8FBF002C,
8FB50028,
8FB40024,
8FB30020,
8FB2001C,
8FB10018,
8FB00014,
03E00008,
27BD0030,
26310001,
00118E00,
00118E03,
A2110044,
1000FFF2,
24020001,
3C040100,
0C400236,
24845334,
1000FFD1,
00000000,
27BDFFE0,
AFB10014,
AFB00010,
AFBF001C,
AFB20018,
00808025,
14800005,
00A08825,
3C040100,
240505FC,
0C400236,
24845334,
16200005,
00000000,
8E020040,
00000000,
14400018,
240505FD,
8E020040,
00000000,
14400004,
240505FE,
3C040100,
0C400236,
24845334,
8E030038,
00000000,
10600007,
00001025,
8E12000C,
02202825,
0C400561,
02002025,
AE12000C,
24020001,
8FBF001C,
8FB20018,
8FB10014,
8FB00010,
03E00008,
27BD0020,
3C040100,
0C400236,
24845334,
1000FFE5,
00000000,
27BDFFE8,
AFB00010,
AFBF0014,
14800005,
00808025,
3C040100,
2405062F,
0C400236,
24845334,
0C400C9C,
00000000,
8E100038,
0C400CAF,
00000000,
8FBF0014,
02001025,
8FB00010,
03E00008,
27BD0018,
27BDFFE0,
AFB10018,
AFBF001C,
AFB00014,
14800005,
00808825,
3C040100,
24050641,
0C400236,
24845334,
0C400C9C,
00000000,
8E220038,
8E30003C,
0C400CAF,
02028023,
8FBF001C,
02001025,
8FB10018,
8FB00014,
03E00008,
27BD0020,
27BDFFE8,
AFB00010,
AFBF0014,
14800005,
00808025,
3C040100,
24050651,
0C400236,
24845334,
8FBF0014,
8E020038,
8FB00010,
03E00008,
27BD0018,
27BDFFE8,
AFB00010,
AFBF0014,
14800005,
00808025,
3C040100,
24050793,
0C400236,
24845334,
8E020038,
8FBF0014,
8FB00010,
2C420001,
03E00008,
27BD0018,
27BDFFE8,
AFB00010,
AFBF0014,
14800005,
00808025,
3C040100,
240507BA,
0C400236,
24845334,
8E030038,
8E02003C,
8FBF0014,
00431026,
8FB00010,
2C420001,
03E00008,
27BD0018,
3C030101,
2463578C,
00001025,
00603025,
2407000A,
8C680000,
00000000,
15000007,
24420001,
2442FFFF,
000210C0,
00C21021,
AC450000,
03E00008,
AC440004,
1447FFF5,
24630008,
03E00008,
00000000,
3C030101,
2463578C,
00001025,
00602825,
2406000A,
8C670004,
00000000,
14E40007,
24420001,
2442FFFF,
000210C0,
00A21021,
8C420000,
03E00008,
00000000,
1446FFF5,
24630008,
03E00008,
00001025,
3C030101,
2463578C,
00001025,
00602825,
2406000A,
8C670004,
00000000,
14E40007,
24420001,
2442FFFF,
000210C0,
00A21021,
AC400000,
03E00008,
AC400004,
1446FFF5,
24630008,
03E00008,
00000000,
27BDFFE8,
AFB00010,
AFBF0014,
14800005,
00808025,
3C040100,
2405065D,
0C400236,
24845334,
0C400968,
02002025,
8FBF0014,
02002025,
8FB00010,
08401323,
27BD0018,
8C820000,
00000000,
10400027,
24870008,
8C820004,
00000000,
8C420004,
00000000,
14470004,
AC820004,
8C82000C,
00000000,
AC820004,
8C820004,
00000000,
8C49000C,
8C820004,
00000000,
8C420004,
00000000,
14E20004,
AC820004,
8C82000C,
00000000,
AC820004,
8C820004,
00A03025,
8C42000C,
00000000,
24430034,
244A0044,
806B0000,
80C80000,
00000000,
150B0005,
00000000,
11000006,
24630001,
146AFFF8,
24C60001,
1522FFE7,
00000000,
00001025,
03E00008,
00000000,
8F828050,
00000000,
8C420000,
00000000,
14400005,
00000000,
2402FFFF,
AF828024,
03E00008,
00000000,
8F828050,
00000000,
8C42000C,
00000000,
8C42000C,
00000000,
8C420004,
1000FFF5,
00000000,
27BDFFE8,
AFB00010,
AFBF0014,
14800005,
00808025,
3C040100,
24050688,
0C400236,
2484534C,
3C030100,
8E040014,
24635450,
14830007,
00001025,
3C030100,
8E040028,
24635478,
10830002,
00000000,
2C820001,
8FBF0014,
8FB00010,
03E00008,
27BD0018,
27BDFFE0,
AFB10014,
AFB00010,
8F918040,
00808025,
8F828018,
8F848018,
AFB20018,
AFBF001C,
24840004,
A0400055,
0C40050E,
00A09025,
2402FFFF,
1602000D,
00000000,
1240000C,
02308021,
8F858018,
8FBF001C,
8FB20018,
8FB10014,
8FB00010,
3C040100,
24A50004,
24845450,
084004E5,
27BD0020,
02308021,
8F828018,
0211882B,
1220000A,
AC500004,
8F84804C,
8F858018,
8FBF001C,
8FB20018,
8FB10014,
8FB00010,
24A50004,
084004F3,
27BD0020,
8F848050,
8F858018,
0C4004F3,
24A50004,
8F828024,
00000000,
0202102B,
10400002,
00000000,
AF908024,
8FBF001C,
8FB20018,
8FB10014,
8FB00010,
03E00008,
27BD0020,
14800003,
00000000,
8F848018,
00000000,
8C82002C,
03E00008,
00000000,
27BDFFE0,
AFB10014,
AFBF001C,
AFB20018,
AFB00010,
14800005,
00808825,
3C040100,
240506E9,
0C400236,
2484534C,
0C4009CB,
02202025,
1040001C,
00008025,
8F82801C,
00000000,
1440001F,
3C040100,
8F828018,
8E30002C,
8C42002C,
26320004,
02402025,
0C40050E,
0202802B,
8E24002C,
8F82803C,
00000000,
0044102B,
10400002,
3A100001,
AF84803C,
00041080,
00441021,
3C040100,
00021080,
248454B4,
02402825,
00822021,
0C4004E5,
00000000,
8FBF001C,
02001025,
8FB20018,
8FB10014,
8FB00010,
03E00008,
27BD0020,
26250018,
1000FFF5,
24845478,
27BDFFE8,
AFBF0014,
0C40024D,
00000000,
8FBF0014,
27BD0018,
AF808038,
08401289,
00000000,
8F82801C,
00000000,
24420001,
AF82801C,
03E00008,
00000000,
8F828040,
03E00008,
00000000,
8F828040,
03E00008,
00000000,
8F828044,
03E00008,
00000000,
27BDFFE8,
AFB00010,
AFBF0014,
14800008,
00808025,
8F908018,
00000000,
16000004,
24050893,
3C040100,
0C400236,
2484534C,
8FBF0014,
26020034,
8FB00010,
03E00008,
27BD0018,
8F828020,
27BDFFE8,
14400005,
AFBF0014,
3C040100,
24050966,
0C400236,
2484534C,
8FBF0014,
8F828020,
03E00008,
27BD0018,
8F82801C,
27BDFFD8,
AFBF0024,
AFB40020,
AFB3001C,
AFB20018,
AFB10014,
1440006D,
AFB00010,
8F918040,
00000000,
26310001,
AF918040,
16200015,
00000000,
8F828050,
00000000,
8C420000,
00000000,
10400004,
240509E4,
3C040100,
0C400236,
2484534C,
8F828050,
8F83804C,
00000000,
AF838050,
AF82804C,
8F82802C,
00000000,
24420001,
AF82802C,
0C4009B8,
00000000,
8F828024,
3C100100,
0222102B,
261054B4,
14400008,
00009825,
8F828050,
00000000,
8C420000,
00000000,
1440001E,
2402FFFF,
AF828024,
8F828018,
00000000,
8C43002C,
00000000,
00031080,
00431021,
00021080,
02028021,
8E020000,
00000000,
2C420002,
14400002,
00000000,
24130001,
8F828030,
00000000,
10400002,
00000000,
24130001,
8FBF0024,
02601025,
8FB40020,
8FB3001C,
8FB20018,
8FB10014,
8FB00010,
03E00008,
27BD0028,
8F828050,
00000000,
8C42000C,
00000000,
8C52000C,
00000000,
8E420004,
00000000,
0222182B,
1460FFD9,
26540004,
0C40050E,
02802025,
8E420028,
00000000,
10400003,
00000000,
0C40050E,
26440018,
8E42002C,
8F83803C,
00000000,
0062182B,
10600002,
00000000,
AF82803C,
00022080,
00822021,
00042080,
02802825,
0C4004E5,
02042021,
8F838018,
8E42002C,
8C63002C,
00000000,
0043102B,
1440FFB7,
00000000,
1000FFB5,
24130001,
8F828034,
00009825,
24420001,
AF828034,
1000FFC4,
00000000,
8F82801C,
27BDFFD8,
AFBF0024,
AFB30020,
AFB2001C,
AFB10018,
1040000A,
AFB00014,
24020001,
AF828030,
8FBF0024,
8FB30020,
8FB2001C,
8FB10018,
8FB00014,
03E00008,
27BD0028,
AF808030,
8F90803C,
3C120100,
00108880,
02308821,
00118880,
265254B4,
3C130100,
02518821,
2673534C,
8E220000,
00000000,
10400018,
00101880,
00701021,
00021080,
02422021,
8C850004,
24420008,
8CA50004,
02421021,
14A20004,
AC850004,
8CA20004,
00000000,
AC820004,
00701821,
00031880,
02439021,
8E420004,
00000000,
8C42000C,
00000000,
AF828018,
AF90803C,
1000FFD5,
00000000,
16000003,
24050B05,
0C400236,
02602025,
2610FFFF,
1000FFDF,
2631FFEC,
27BDFFE0,
AFB10018,
AFB00014,
AFBF001C,
00808025,
14800005,
00A08825,
3C040100,
24050B15,
0C400236,
2484534C,
8F858018,
02002025,
0C4004F3,
24A50018,
8FBF001C,
8FB00014,
02202025,
8FB10018,
24050001,
084009E3,
27BD0020,
27BDFFE0,
AFB20018,
AFB10014,
AFB00010,
AFBF001C,
00808825,
00A08025,
14800005,
00C09025,
3C040100,
24050B26,
0C400236,
2484534C,
8F82801C,
00000000,
14400004,
3C040100,
24050B2A,
0C400236,
2484534C,
8F828018,
3C038000,
8F858018,
02038025,
02202025,
AC500018,
0C4004E5,
24A50018,
8FBF001C,
8FB10014,
8FB00010,
02402025,
8FB20018,
24050001,
084009E3,
27BD0020,
8C82000C,
27BDFFE0,
AFB00014,
8C50000C,
AFBF001C,
16000005,
AFB10018,
3C040100,
24050B70,
0C400236,
2484534C,
26110018,
0C40050E,
02202025,
8F82801C,
00000000,
14400022,
3C040100,
26110004,
0C40050E,
02202025,
8E04002C,
8F82803C,
00000000,
0044102B,
10400002,
00000000,
AF84803C,
00041080,
00441021,
3C040100,
00021080,
248454B4,
02202825,
00822021,
0C4004E5,
00000000,
8F828018,
8E03002C,
8C42002C,
00000000,
0043182B,
10600003,
00001025,
24020001,
AF828030,
8FBF001C,
8FB10018,
8FB00014,
03E00008,
27BD0020,
02202825,
1000FFEE,
24845478,
8F82801C,
27BDFFE0,
AFB10018,
AFB00014,
AFBF001C,
00808825,
14400005,
00A08025,
3C040100,
24050BA8,
0C400236,
2484534C,
3C028000,
02028025,
AE300000,
8E30000C,
00000000,
16000004,
24050BB0,
3C040100,
0C400236,
2484534C,
02202025,
0C40050E,
26110004,
0C40050E,
02202025,
8E04002C,
8F82803C,
00000000,
0044102B,
10400002,
00000000,
AF84803C,
00041080,
00441021,
3C040100,
00021080,
248454B4,
00822021,
0C4004E5,
02202825,
8F828018,
8E03002C,
8C42002C,
00000000,
0043182B,
10600003,
00001025,
24020001,
AF828030,
8FBF001C,
8FB10018,
8FB00014,
03E00008,
27BD0020,
27BDFFE8,
AFB00010,
AFBF0014,
14800005,
00808025,
3C040100,
24050BD0,
0C400236,
2484534C,
8F82802C,
8FBF0014,
AE020000,
8F828040,
00000000,
AE020004,
8FB00010,
03E00008,
27BD0018,
24020001,
AF828030,
03E00008,
00000000,
14800003,
00000000,
8F848018,
00000000,
8C840030,
240500A5,
00801825,
90660000,
00000000,
10C50004,
00641023,
00021082,
03E00008,
3042FFFF,
1000FFF8,
24630001,
8F828018,
03E00008,
00000000,
8F838038,
00000000,
10600005,
24020001,
8F82801C,
00000000,
2C420001,
00021040,
03E00008,
00000000,
1080003E,
00000000,
8F828018,
8C83002C,
8C42002C,
27BDFFE0,
0062102B,
AFBF001C,
AFB20018,
AFB10014,
1040002F,
AFB00010,
8C820018,
00000000,
04400008,
00031080,
8F828018,
00000000,
8C45002C,
24020005,
00451023,
AC820018,
00031080,
00431021,
3C110100,
00021080,
263154B4,
8C830014,
02221021,
14620017,
24920004,
00808025,
0C40050E,
02402025,
8F828018,
8F83803C,
8C42002C,
00000000,
0062182B,
10600002,
AE02002C,
AF82803C,
00022080,
00822021,
00042080,
8FBF001C,
8FB00010,
02402825,
02242021,
8FB20018,
8FB10014,
084004E5,
27BD0020,
8F828018,
00000000,
8C42002C,
00000000,
AC82002C,
8FBF001C,
8FB20018,
8FB10014,
8FB00010,
27BD0020,
03E00008,
00000000,
14800009,
00001025,
03E00008,
00000000,
00001025,
8FBF001C,
8FB10018,
8FB00014,
03E00008,
27BD0020,
8F828018,
27BDFFE0,
AFB00014,
AFBF001C,
AFB10018,
10820005,
00808025,
3C040100,
24050ED6,
0C400236,
2484534C,
8E02004C,
00000000,
14400005,
3C040100,
24050ED8,
0C400236,
2484534C,
8E02004C,
8E04002C,
8E030048,
2442FFFF,
1083FFE3,
AE02004C,
1440FFE2,
00001025,
26110004,
0C40050E,
02202025,
8E040048,
24020005,
00441023,
AE020018,
8F82803C,
00000000,
0044102B,
10400002,
AE04002C,
AF84803C,
00041080,
00442021,
3C020100,
244254B4,
00042080,
00442021,
0C4004E5,
02202825,
1000FFCB,
24020001,
27BDFFE8,
AFBF0014,
0C40024D,
00000000,
8F828038,
00000000,
10400008,
00000000,
8F838018,
00000000,
8C620044,
00000000,
24420001,
AC620044,
8F828018,
8FBF0014,
00000000,
03E00008,
27BD0018,
8F828038,
00000000,
10400015,
00000000,
8F828018,
00000000,
8C420044,
00000000,
1040000F,
00000000,
8F838018,
00000000,
8C620044,
00000000,
2442FFFF,
AC620044,
8F828018,
00000000,
8C420044,
00000000,
14400003,
00000000,
08400248,
00000000,
03E00008,
00000000,
27BDFFC8,
AFB2001C,
00069080,
AFB40024,
0080A025,
02402025,
AFB70030,
AFB50028,
AFB30020,
AFB10018,
AFBF0034,
AFB6002C,
AFB00014,
00A08825,
8FB3004C,
0C4012B1,
00E0A825,
1040008F,
2417FFFF,
24040058,
0C4012B1,
0040B025,
10400087,
00408025,
02403025,
240500A5,
AC560030,
0C401438,
02C02025,
2642FFFC,
8E120030,
02202825,
02429021,
2402FFFC,
02429024,
26230010,
26020034,
80A40000,
00000000,
A0440000,
80A40000,
00000000,
10800003,
24A50001,
1465FFF8,
24420001,
8FB60048,
00000000,
2EC20005,
14400002,
A2000043,
24160004,
26110004,
AE16002C,
AE160048,
02202025,
0C4004E3,
AE00004C,
0C4004E3,
26040018,
24020005,
0056B023,
AE000050,
AE100010,
AE160018,
AE100024,
AE000044,
A2000054,
A2000055,
02A03025,
02802825,
0C400085,
02402025,
12600002,
AE020000,
AE700000,
0C400C9C,
00000000,
8F828044,
3C120100,
24420001,
AF828044,
8F828018,
00000000,
14400058,
00000000,
AF908018,
8F838044,
24020001,
14620022,
00000000,
0C4004DB,
264454B4,
3C040100,
0C4004DB,
248454C8,
3C040100,
0C4004DB,
248454DC,
3C040100,
0C4004DB,
248454F0,
3C040100,
24845504,
0C4004DB,
3C140100,
3C130100,
0C4004DB,
268454A0,
0C4004DB,
2664548C,
3C040100,
0C4004DB,
24845478,
3C040100,
0C4004DB,
24845464,
3C040100,
24845450,
269454A0,
0C4004DB,
2673548C,
AF948050,
AF93804C,
8F828028,
8E04002C,
24420001,
AF828028,
8F82803C,
00000000,
0044102B,
10400003,
00041080,
AF84803C,
00041080,
00441021,
00021080,
264454B4,
00822021,
0C4004E5,
02202825,
0C400CAF,
00000000,
8F828038,
00000000,
1040000F,
24170001,
8F828018,
8E03002C,
8C42002C,
00000000,
0043102B,
10400008,
00000000,
0C400120,
00000000,
10000004,
00000000,
0C401323,
02C02025,
2417FFFF,
8FBF0034,
02E01025,
8FB6002C,
8FB70030,
8FB50028,
8FB40024,
8FB30020,
8FB2001C,
8FB10018,
8FB00014,
03E00008,
27BD0038,
8F828038,
00000000,
1440FFCC,
00000000,
8F828018,
8E03002C,
8C42002C,
00000000,
0062102B,
1440FFC5,
00000000,
AF908018,
1000FFC2,
00000000,
27BDFFE0,
27828020,
3C050100,
3C040100,
00003825,
AFA20014,
AFA00010,
2406012C,
24A55364,
AFB00018,
AFBF001C,
0C400CC9,
24844008,
00408025,
24020001,
1602000C,
2402FFFF,
0C40024D,
00000000,
2402FFFF,
AF828024,
8FBF001C,
AF908038,
8FB00018,
27BD0020,
AF808040,
0840127D,
00000000,
16020007,
3C040100,
8FBF001C,
8FB00018,
2405078B,
2484534C,
08400236,
27BD0020,
8FBF001C,
8FB00018,
03E00008,
27BD0020,
27BDFFE0,
AFB00014,
00808025,
AFBF001C,
0C400C9C,
AFB10018,
16000004,
26110004,
8F908018,
00000000,
26110004,
0C40050E,
02202025,
8E020028,
00000000,
10400003,
00000000,
0C40050E,
26040018,
8F828028,
00000000,
24420001,
AF828028,
8F828018,
00000000,
1602001E,
02202825,
3C040100,
0C4004E5,
24845464,
8F828048,
00000000,
24420001,
AF828048,
0C400CAF,
00000000,
8F828038,
00000000,
1040001D,
00000000,
8F828018,
00000000,
16020019,
00000000,
8F82801C,
00000000,
10400004,
24050465,
3C040100,
0C400236,
2484534C,
8FBF001C,
8FB10018,
8FB00014,
08400120,
27BD0020,
8F828044,
8E040030,
2442FFFF,
AF828044,
0C401323,
00000000,
0C401323,
02002025,
0C4009B8,
00000000,
1000FFDF,
00000000,
8FBF001C,
8FB10018,
8FB00014,
03E00008,
27BD0020,
27BDFFE0,
AFB10018,
AFBF001C,
AFB00014,
14800005,
00808825,
3C040100,
24050502,
0C400236,
2484534C,
8F838018,
00000000,
12230016,
00001025,
0C400C9C,
00000000,
8E300014,
0C400CAF,
00000000,
8F838050,
00000000,
1203000D,
24020002,
8F83804C,
00000000,
12030009,
00000000,
3C020100,
24425450,
1602000A,
3C030100,
8E220028,
00000000,
2C420001,
24420002,
8FBF001C,
8FB10018,
8FB00014,
03E00008,
27BD0020,
24635464,
1203FFF9,
24020004,
1200FFF7,
00000000,
1000FFF5,
24020001,
27BDFFE8,
AFB00010,
AFBF0014,
0C400C9C,
00808025,
16000003,
02002025,
8F848018,
00000000,
8C90002C,
0C400CAF,
00000000,
8FBF0014,
02001025,
8FB00010,
03E00008,
27BD0018,
27BDFFD8,
2CA20005,
AFB2001C,
AFB00014,
AFBF0024,
AFB30020,
AFB10018,
00808025,
14400006,
00A09025,
3C040100,
24050587,
0C400236,
2484534C,
24120004,
0C400C9C,
00000000,
16000003,
00000000,
8F908018,
00000000,
8E020048,
00000000,
12420035,
0052182B,
1060003A,
00000000,
8F838018,
00000000,
12030007,
00008825,
8F838018,
00000000,
8C71002C,
00000000,
0251882B,
3A310001,
8E03002C,
00000000,
14430002,
00000000,
AE12002C,
8E020018,
00000000,
04400004,
AE120048,
24050005,
00B29023,
AE120018,
00031080,
00431021,
3C120100,
00021080,
265254B4,
8E030014,
02421021,
14620010,
26130004,
0C40050E,
02602025,
8E02002C,
8F83803C,
00000000,
0062182B,
10600002,
00000000,
AF82803C,
00022080,
00822021,
00042080,
02602825,
0C4004E5,
02442021,
12200003,
00000000,
0C400120,
00000000,
8FBF0024,
8FB30020,
8FB2001C,
8FB10018,
8FB00014,
08400CAF,
27BD0028,
8F918018,
00000000,
02118826,
1000FFCD,
2E310001,
27BDFFE0,
AFB00014,
00808025,
AFBF001C,
0C400C9C,
AFB10018,
16000004,
26110004,
8F908018,
00000000,
26110004,
0C40050E,
02202025,
8E020028,
00000000,
10400004,
02202825,
0C40050E,
26040018,
02202825,
3C110100,
0C4004E5,
26245450,
0C400CAF,
00000000,
8F828038,
00000000,
10400007,
00000000,
0C400C9C,
00000000,
0C4009B8,
00000000,
0C400CAF,
00000000,
8F828018,
00000000,
16020017,
00000000,
8F828038,
00000000,
1040000D,
00000000,
8F82801C,
00000000,
10400004,
3C040100,
2405065E,
0C400236,
2484534C,
8FBF001C,
8FB10018,
8FB00014,
08400120,
27BD0020,
8F828044,
8E235450,
00000000,
14620007,
00000000,
AF808018,
8FBF001C,
8FB10018,
8FB00014,
03E00008,
27BD0020,
8FBF001C,
8FB10018,
8FB00014,
08400B08,
27BD0020,
14800029,
240506B2,
3C040100,
08400236,
2484534C,
0C400C9C,
00808025,
0C4009CB,
02002025,
1040001B,
26110004,
0C40050E,
02202025,
8E04002C,
8F82803C,
00000000,
0044102B,
10400003,
00041080,
AF84803C,
00041080,
00441021,
3C040100,
00021080,
248454B4,
00822021,
0C4004E5,
02202825,
8F838018,
8E02002C,
8C63002C,
00000000,
0043102B,
14400003,
00000000,
0C400120,
00000000,
8FBF001C,
8FB10018,
8FB00014,
08400CAF,
27BD0020,
8F828018,
27BDFFE0,
AFBF001C,
AFB10018,
1482FFD6,
AFB00014,
8FBF001C,
8FB10018,
8FB00014,
03E00008,
27BD0020,
8F82801C,
27BDFFD0,
AFBF002C,
AFB50028,
AFB40024,
AFB30020,
AFB2001C,
AFB10018,
14400005,
AFB00014,
3C040100,
240507EF,
0C400236,
2484534C,
0C400C9C,
00000000,
8F82801C,
00000000,
2442FFFF,
AF82801C,
8F82801C,
00000000,
1040000E,
00000000,
00008025,
0C400CAF,
00000000,
8FBF002C,
02001025,
8FB50028,
8FB40024,
8FB30020,
8FB2001C,
8FB10018,
8FB00014,
03E00008,
27BD0030,
8F828044,
00000000,
1040FFF0,
3C140100,
3C110100,
00008025,
26925478,
263154B4,
24130001,
8E825478,
00000000,
1440001A,
00000000,
12000003,
00000000,
0C4009B8,
00000000,
8F908034,
00000000,
1200000A,
24110001,
0C400A8D,
00000000,
10400002,
00000000,
AF918030,
2610FFFF,
1600FFF9,
00000000,
AF808034,
8F828030,
00000000,
1040FFD2,
00000000,
0C400120,
24100001,
1000FFCF,
00000000,
8E42000C,
00000000,
8C50000C,
00000000,
26040018,
0C40050E,
26150004,
0C40050E,
02A02025,
8E02002C,
8F83803C,
00000000,
0062182B,
10600002,
00000000,
AF82803C,
00022080,
00822021,
00042080,
02A02825,
0C4004E5,
02242021,
8F838018,
8E02002C,
8C63002C,
00000000,
0043102B,
1440FFC7,
00000000,
AF938030,
1000FFC4,
00000000,
27BDFFE0,
AFB10018,
AFB00014,
AFBF001C,
00808825,
14800005,
00A08025,
3C040100,
24050479,
0C400236,
2484534C,
16000004,
2405047A,
3C040100,
0C400236,
2484534C,
8F82801C,
00000000,
10400004,
3C040100,
2405047B,
0C400236,
2484534C,
0C400A61,
00000000,
8E230000,
8F848040,
02038021,
0083282B,
10A00005,
0203182B,
10600005,
00002825,
10000003,
0090282B,
1060FFFD,
24050001,
10A00004,
AE300000,
00002825,
0C4009E3,
02042023,
0C400F0A,
00000000,
14400006,
00000000,
8FBF001C,
8FB10018,
8FB00014,
08400120,
27BD0020,
8FBF001C,
8FB10018,
8FB00014,
03E00008,
27BD0020,
14800007,
00000000,
08400120,
00000000,
8FBF0014,
8FB00010,
1000FFFB,
27BD0018,
8F82801C,
27BDFFE8,
AFB00010,
AFBF0014,
10400005,
00808025,
3C040100,
240504D6,
0C400236,
2484534C,
0C400A61,
00002825,
0C4009E3,
02002025,
0C400F0A,
00000000,
1040FFEB,
00000000,
8FBF0014,
8FB00010,
03E00008,
27BD0018,
27BDFFE0,
AFB10018,
AFBF001C,
AFB00014,
0C40147F,
00808825,
2C420010,
14400004,
240508DD,
3C040100,
0C400236,
2484534C,
0C400A61,
3C0D0100,
00006025,
25AD54B4,
240EFF9C,
25840050,
02202825,
0C40098B,
01A42021,
14400019,
00408025,
258CFFEC,
158EFFF9,
25840050,
8F848050,
0C40098B,
02202825,
14400011,
00408025,
8F84804C,
0C40098B,
02202825,
1440000C,
00408025,
3C040100,
02202825,
0C40098B,
24845450,
14400006,
00408025,
3C040100,
02202825,
0C40098B,
24845464,
00408025,
0C400F0A,
00000000,
8FBF001C,
02001025,
8FB10018,
8FB00014,
03E00008,
27BD0020,
27BDFFD8,
AFB10018,
3C110100,
AFB30020,
AFB2001C,
AFBF0024,
AFB00014,
26335464,
3C120100,
8F828048,
00000000,
1440000A,
00000000,
8E4254B4,
00000000,
2C420002,
1440FFF8,
00000000,
0C400120,
00000000,
1000FFF4,
00000000,
0C400A61,
00000000,
8E305464,
0C400F0A,
00000000,
1200FFED,
00000000,
0C400C9C,
00000000,
8E62000C,
00000000,
8C50000C,
0C40050E,
26040004,
8F828044,
00000000,
2442FFFF,
AF828044,
8F828048,
00000000,
2442FFFF,
AF828048,
0C400CAF,
00000000,
8E040030,
0C401323,
00000000,
0C401323,
02002025,
1000FFD5,
00000000,
27BDFFE0,
AFB00014,
AFBF001C,
AFB10018,
14800005,
00808025,
3C040100,
24050987,
0C400236,
2484534C,
0C400A61,
02002025,
0C400DF5,
00000000,
24030002,
14430026,
26110004,
0C40050E,
02202025,
0C400C9C,
00000000,
8E020028,
00000000,
10400005,
00000000,
0C40050E,
26040018,
24020001,
A2020055,
0C400CAF,
00000000,
8E04002C,
8F82803C,
00000000,
0044102B,
10400003,
00041080,
AF84803C,
00041080,
00441021,
3C040100,
00021080,
248454B4,
00822021,
0C4004E5,
02202825,
8F838018,
8E02002C,
8C63002C,
00000000,
0062102B,
10400002,
24020001,
AF828030,
0C400F0A,
00000000,
8FBF001C,
8FB10018,
8FB00014,
00001025,
03E00008,
27BD0020,
27BDFFE0,
AFB20018,
AFB10014,
AFBF001C,
AFB00010,
00808825,
14800005,
00A09025,
3C040100,
24050BDA,
0C400236,
2484534C,
16400004,
3C040100,
24050BDB,
0C400236,
2484534C,
0C400C9C,
00000000,
8F848040,
8F828018,
00000000,
90420055,
00000000,
1040000D,
2402FFFF,
8F828018,
24100001,
A0400055,
0C400CAF,
00000000,
8FBF001C,
02001025,
8FB20018,
8FB10014,
8FB00010,
03E00008,
27BD0020,
8E430000,
00000000,
1062FFF4,
00008025,
8F85802C,
8E260000,
8E220004,
10C50003,
0082282B,
10A0FFED,
24100001,
00822823,
00A3282B,
10A0FFE9,
24100001,
00641823,
00621821,
AE430000,
0C400BED,
02202025,
1000FFE2,
00008025,
8F828018,
8F848018,
8F838018,
8C420018,
8C65002C,
24030005,
00651823,
03E00008,
AC830018,
8F828018,
00000000,
10400007,
00000000,
8F838018,
00000000,
8C62004C,
00000000,
24420001,
AC62004C,
8F828018,
03E00008,
00000000,
27BDFFE0,
AFB10018,
AFB00014,
AFBF001C,
00808825,
0C400C9C,
00A08025,
8F828018,
00000000,
8C420050,
00000000,
1440000A,
00000000,
8F828018,
24030001,
A0430054,
12000005,
24050001,
0C4009E3,
02002025,
0C400120,
00000000,
0C400CAF,
00000000,
0C400C9C,
00000000,
8F828018,
00000000,
8C500050,
00000000,
12000005,
00000000,
8F828018,
1220000D,
2603FFFF,
AC400050,
8F828018,
00000000,
A0400054,
0C400CAF,
00000000,
8FBF001C,
02001025,
8FB10018,
8FB00014,
03E00008,
27BD0020,
AC430050,
1000FFF3,
00000000,
27BDFFD8,
AFB30020,
AFB2001C,
AFB10018,
AFB00014,
AFBF0024,
00808825,
00A08025,
00C09025,
0C400C9C,
00E09825,
8F828018,
24030002,
90420054,
00000000,
304200FF,
10430010,
00000000,
8F828018,
00118827,
8C440050,
24030001,
02248824,
AC510050,
8F828018,
00000000,
A0430054,
12600005,
24050001,
0C4009E3,
02602025,
0C400120,
00000000,
0C400CAF,
00000000,
0C400C9C,
00000000,
12400006,
00000000,
8F828018,
00000000,
8C420050,
00000000,
AE420000,
8F828018,
00008825,
90430054,
24020001,
306300FF,
10620007,
00000000,
8F828018,
00108027,
8C430050,
24110001,
02038024,
AC500050,
8F828018,
00000000,
A0400054,
0C400CAF,
00000000,
8FBF0024,
02201025,
8FB30020,
8FB2001C,
8FB10018,
8FB00014,
03E00008,
27BD0028,
27BDFFD8,
AFB30020,
AFB2001C,
AFB10018,
AFB00014,
AFBF0024,
00808025,
00A09025,
00C08825,
14800005,
00E09825,
3C040100,
2405110C,
0C400236,
2484534C,
0C400C9C,
00000000,
12600004,
00000000,
8E020050,
00000000,
AE620000,
92030054,
24020002,
A2020054,
24020002,
12220023,
306300FF,
2E240003,
10800009,
00000000,
24020001,
12220017,
00000000,
24020001,
10620020,
00000000,
10000008,
24110001,
24040003,
12240012,
24040004,
1624FFF7,
00000000,
1462000E,
00008825,
0C400CAF,
00000000,
8FBF0024,
02201025,
8FB30020,
8FB2001C,
8FB10018,
8FB00014,
03E00008,
27BD0028,
8E020050,
00000000,
00529025,
AE120050,
1000FFE6,
24020001,
8E020050,
00000000,
24420001,
AE020050,
1000FFE0,
24020001,
26110004,
0C40050E,
02202025,
8E04002C,
8F82803C,
00000000,
0044102B,
10400003,
00041080,
AF84803C,
00041080,
00441021,
3C040100,
00021080,
248454B4,
00822021,
0C4004E5,
02202825,
8E020028,
00000000,
10400004,
3C040100,
24051144,
0C400236,
2484534C,
8F838018,
8E02002C,
8C63002C,
00000000,
0062102B,
1040FFC2,
00000000,
0C400120,
24110001,
1000FFC7,
00000000,
27BDFFD8,
AFB40020,
AFB3001C,
AFB20018,
AFB10014,
AFB00010,
AFBF0024,
00808025,
00A09825,
00C08825,
8FB20038,
14800005,
00E0A025,
3C040100,
24051177,
0C400236,
2484534C,
12800004,
00000000,
8E020050,
00000000,
AE820000,
92030054,
24020002,
24040002,
306300FF,
A2020054,
12240021,
00000000,
2E220003,
10400009,
24020003,
24020001,
12220015,
00000000,
24020001,
1062001E,
00000000,
10000008,
24020001,
12220011,
00000000,
24020004,
1622FFF7,
00000000,
1464000C,
00001025,
8FBF0024,
8FB40020,
8FB3001C,
8FB20018,
8FB10014,
8FB00010,
03E00008,
27BD0028,
8E020050,
00000000,
00539825,
AE130050,
1000FFE8,
24020001,
8E020050,
00000000,
24420001,
AE020050,
1000FFE2,
24020001,
8E020028,
00000000,
10400004,
240511BE,
3C040100,
0C400236,
2484534C,
8F82801C,
00000000,
1440001F,
3C040100,
26110004,
0C40050E,
02202025,
8E04002C,
8F82803C,
00000000,
0044102B,
10400003,
00041080,
AF84803C,
00041080,
00441021,
3C040100,
00021080,
248454B4,
02202825,
00822021,
0C4004E5,
00000000,
8F838018,
8E02002C,
8C63002C,
00000000,
0062102B,
1040FFBF,
00000000,
12400006,
24020001,
1000FFC4,
AE420000,
26050018,
1000FFF1,
24845478,
AF828030,
1000FFBE,
00000000,
27BDFFE0,
AFB10014,
AFB00010,
AFBF001C,
AFB20018,
00808025,
14800005,
00A08825,
3C040100,
240511F2,
0C400236,
2484534C,
24030002,
92020054,
A2030054,
8E030050,
304200FF,
24630001,
AE030050,
24030001,
14430029,
00000000,
8E020028,
00000000,
10400004,
24051218,
3C040100,
0C400236,
2484534C,
8F82801C,
00000000,
14400024,
3C040100,
26120004,
0C40050E,
02402025,
8E04002C,
8F82803C,
00000000,
0044102B,
10400003,
00041080,
AF84803C,
00041080,
00441021,
3C040100,
00021080,
248454B4,
02402825,
00822021,
0C4004E5,
00000000,
8F838018,
8E02002C,
8C63002C,
00000000,
0062102B,
10400004,
00000000,
1220000B,
24020001,
AE220000,
8FBF001C,
8FB20018,
8FB10014,
8FB00010,
03E00008,
27BD0020,
26050018,
1000FFEC,
24845478,
AF828030,
1000FFF5,
00000000,
27BDFFE0,
AFB00014,
AFBF001C,
AFB10018,
14800002,
00808025,
8F908018,
0C400C9C,
00000000,
92030054,
24020002,
306300FF,
14620003,
00008825,
A2000054,
24110001,
0C400CAF,
00000000,
8FBF001C,
02201025,
8FB00014,
8FB10018,
03E00008,
27BD0020,
03E00008,
00000000,
27BDFFE8,
AFBF0014,
0C4000E7,
00000000,
0C400248,
00000000,
0C4000F6,
00000000,
0C40024D,
00000000,
1000FFFF,
00000000,
3C040100,
24050070,
08400236,
2484536C,
27828068,
8C430000,
00000000,
0064282B,
14A0001D,
00000000,
8C450004,
00000000,
00453021,
14860006,
00000000,
8C840004,
00000000,
00852021,
AC440004,
00402025,
8C860004,
00000000,
00862821,
14650009,
00000000,
8F858064,
00000000,
10650005,
00000000,
8C650004,
8C630000,
00A62821,
AC850004,
10820002,
AC830000,
AC440000,
03E00008,
00000000,
1000FFDE,
00601025,
27BDFFD8,
AFB00014,
AFBF0024,
AFB30020,
AFB2001C,
AFB10018,
0C400A61,
00808025,
8F828064,
00000000,
14400012,
3C050100,
24A35518,
3402FFF8,
2404FFFC,
00621021,
00441024,
00432023,
AF80806C,
AF838068,
AC400004,
AC400000,
AF828064,
ACA25518,
3C028000,
AC640004,
AF84805C,
AF848060,
AF828058,
8F828058,
00000000,
02021024,
1440003A,
00009025,
12000038,
26100008,
32020003,
10400003,
2404FFFC,
02048024,
26100004,
12000031,
00009025,
8F828060,
00000000,
0050102B,
1440002C,
27838068,
8F918068,
00000000,
8E220004,
00000000,
0050202B,
14800035,
00000000,
8F848064,
00000000,
12240021,
00009025,
8C720000,
8E240000,
00501023,
2C420011,
26520008,
1440000E,
AC640000,
02309821,
32620003,
10400004,
3C040100,
240500EC,
0C400236,
24845384,
8E220004,
02602025,
00501023,
AE620004,
0C40128D,
AE300004,
8F828060,
8E240004,
8F83805C,
00441023,
0043182B,
10600002,
AF828060,
AF82805C,
8F828058,
AE200000,
00441025,
AE220004,
0C400F0A,
00000000,
32420003,
10400004,
2405012C,
3C040100,
0C400236,
24845384,
8FBF0024,
02401025,
8FB30020,
8FB2001C,
8FB10018,
8FB00014,
03E00008,
27BD0028,
8E240000,
00000000,
1080FFC9,
00000000,
02201825,
1000FFC1,
00808825,
1080002E,
00000000,
8C82FFFC,
8F838058,
27BDFFE8,
00431024,
AFB00010,
AFBF0014,
14400005,
00808025,
3C040100,
24050140,
0C400236,
24845384,
8E02FFF8,
00000000,
10400004,
3C040100,
24050141,
0C400236,
24845384,
8E03FFFC,
8F828058,
00000000,
00622024,
10800012,
00000000,
8E04FFF8,
00000000,
1480000E,
00021027,
00431024,
0C400A61,
AE02FFFC,
8E03FFFC,
8F828060,
2604FFF8,
00431021,
0C40128D,
AF828060,
8FBF0014,
8FB00010,
08400F0A,
27BD0018,
8FBF0014,
8FB00010,
27BD0018,
03E00008,
00000000,
8F828060,
03E00008,
00000000,
8F82805C,
03E00008,
00000000,
03E00008,
00000000,
28CA0008,
1540005B,
00801025,
00A4C026,
33180003,
17000066,
00043823,
30E70003,
10E00005,
00C73023,
88B80000,
00A72821,
A8980000,
00872021,
30D8003F,
10D80026,
00D83823,
00873821,
8CA80000,
8CA90004,
8CAA0008,
8CAB000C,
8CAC0010,
8CAD0014,
8CAE0018,
8CAF001C,
AC880000,
AC890004,
AC8A0008,
AC8B000C,
AC8C0010,
AC8D0014,
AC8E0018,
AC8F001C,
8CA80020,
8CA90024,
8CAA0028,
8CAB002C,
8CAC0030,
8CAD0034,
8CAE0038,
8CAF003C,
AC880020,
AC890024,
AC8A0028,
AC8B002C,
AC8C0030,
AC8D0034,
AC8E0038,
AC8F003C,
24840040,
1487FFDE,
24A50040,
03003025,
30D8001F,
10D80013,
00000000,
8CA80000,
8CA90004,
8CAA0008,
8CAB000C,
8CAC0010,
8CAD0014,
8CAE0018,
8CAF001C,
24A50020,
AC880000,
AC890004,
AC8A0008,
AC8B000C,
AC8C0010,
AC8D0014,
AC8E0018,
AC8F001C,
24840020,
33060003,
10D80007,
03063823,
00873821,
8CAB0000,
24840004,
24A50004,
1487FFFC,
AC8BFFFC,
18C00006,
00863821,
80A30000,
24840001,
24A50001,
1487FFFC,
A083FFFF,
03E00008,
00000000,
30D80003,
1306FFF5,
30990003,
1720FFF3,
30B90003,
1720FFF1,
00D83823,
00873821,
8CAB0000,
24840004,
24A50004,
1487FFFC,
AC8BFFFC,
1000FFE9,
03003025,
30E70003,
10E00006,
00C73023,
88A30000,
98A30003,
00A72821,
A8830000,
00872021,
30D8003F,
10D80036,
00D83823,
00873821,
88A80000,
88A90004,
88AA0008,
88AB000C,
88AC0010,
88AD0014,
88AE0018,
88AF001C,
98A80003,
98A90007,
98AA000B,
98AB000F,
98AC0013,
98AD0017,
98AE001B,
98AF001F,
AC880000,
AC890004,
AC8A0008,
AC8B000C,
AC8C0010,
AC8D0014,
AC8E0018,
AC8F001C,
88A80020,
88A90024,
88AA0028,
88AB002C,
88AC0030,
88AD0034,
88AE0038,
88AF003C,
98A80023,
98A90027,
98AA002B,
98AB002F,
98AC0033,
98AD0037,
98AE003B,
98AF003F,
AC880020,
AC890024,
AC8A0028,
AC8B002C,
AC8C0030,
AC8D0034,
AC8E0038,
AC8F003C,
24840040,
1487FFCE,
24A50040,
03003025,
30D8001F,
10D8001B,
00000000,
88A80000,
88A90004,
88AA0008,
88AB000C,
88AC0010,
88AD0014,
88AE0018,
88AF001C,
98A80003,
98A90007,
98AA000B,
98AB000F,
98AC0013,
98AD0017,
98AE001B,
98AF001F,
24A50020,
AC880000,
AC890004,
AC8A0008,
AC8B000C,
AC8C0010,
AC8D0014,
AC8E0018,
AC8F001C,
24840020,
33060003,
10D80008,
03063823,
00873821,
88A30000,
98A30003,
24840004,
24A50004,
1487FFFB,
AC83FFFC,
10C0FF87,
00863821,
80A30000,
24840001,
24A50001,
1487FFFC,
A083FFFF,
03E00008,
00000000,
28CA0008,
1540003E,
00801025,
10A00007,
00043823,
00000000,
30A500FF,
00055200,
00AA2825,
00055400,
00AA2825,
30EA0003,
11400003,
00CA3023,
A8850000,
008A2021,
30EA0004,
11400003,
00CA3023,
AC850000,
008A2021,
30D8003F,
10D80016,
00D83823,
00873821,
AC850000,
AC850004,
AC850008,
AC85000C,
AC850010,
AC850014,
AC850018,
AC85001C,
AC850020,
AC850024,
AC850028,
AC85002C,
AC850030,
AC850034,
AC850038,
AC85003C,
24840040,
1487FFEE,
00000000,
03003025,
30D8001F,
10D8000A,
00000000,
AC850000,
AC850004,
AC850008,
AC85000C,
AC850010,
AC850014,
AC850018,
AC85001C,
24840020,
33060003,
10D80005,
03063823,
00873821,
24840004,
1487FFFE,
AC85FFFC,
18C00004,
00863821,
24840001,
1487FFFE,
A085FFFF,
03E00008,
00000000,
24820001,
90830000,
00000000,
1460FFFD,
24840001,
03E00008,
00821023,
2A2A2A2A,
20546872,
6561642D,
4D657472,
69632050,
7265656D,
70746976,
65205363,
68656475,
6C696E67,
20546573,
74202A2A,
2A2A2052,
656C6174,
69766520,
54696D65,
3A202575,
0A0D0000,
4552524F,
523A2049,
6E76616C,
69642063,
6F756E74,
65722076,
616C7565,
2873292E,
20507265,
656D7074,
69766520,
636F756E,
74657273,
2073686F,
756C6420,
6E6F7420,
6265206D,
6F726520,
74686174,
20312064,
69666665,
72656E74,
20746861,
6E207468,
65206176,
65726167,
65210A0D,
00000000,
54696D65,
20506572,
696F6420,
546F7461,
6C3A2020,
25750A0D,
0A0D0000,
416C6976,
652E2E2E,
0A0D0000,
41737365,
72743A0A,
0D4D6573,
73616765,
3A25730A,
0D4C696E,
653A2564,
0A0D0000,
746D5F70,
6F727469,
6E675F6C,
61796572,
5F667265,
6572746F,
732E6300,
2E2E2F2E,
2E2F6672,
65657274,
6F732F71,
75657565,
2E630000,
2E2E2F2E,
2E2F6672,
65657274,
6F732F74,
61736B73,
2E630000,
49444C45,
00000000,
2E2E2F2E,
2E2F6672,
65657274,
6F732F70,
6F72742E,
63000000,
2E2E2F2E,
2E2F6672,
65657274,
6F732F68,
6561705F,
342E6300,
00000000,
00000100,
01010001,
00000000,
00000000,
00000000,
00000000;
