----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 02/14/2017 02:57:27 PM
-- Design Name: 
-- Module Name: plasoc_axi4_full2lite_pack - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

package plasoc_axi4_full2lite_pack is

    constant axi_burst_fixed : std_logic_vector := "00";
    constant axi_burst_incr : std_logic_vector := "01";
    
end package;