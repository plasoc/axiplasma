library ieee;
use ieee.std_logic_1164.all;

package bram_pack is

	constant cpu_width : integer := 32;
	constant ram_size : integer := 16384;
	subtype word_type is std_logic_vector(cpu_width-1 downto 0);
	type ram_type is array(0 to ram_size-1) of word_type;
	function load_hex return ram_type;

end package;

package body bram_pack is

	function load_hex return ram_type is
		variable ram_buffer : ram_type := (others=>(others=>'0'));
	begin
		ram_buffer(0) := X"3C1C0101";
		ram_buffer(1) := X"279C8830";
		ram_buffer(2) := X"3C050100";
		ram_buffer(3) := X"24A50840";
		ram_buffer(4) := X"3C040100";
		ram_buffer(5) := X"24840A94";
		ram_buffer(6) := X"3C1D0100";
		ram_buffer(7) := X"27BD0A38";
		ram_buffer(8) := X"ACA00000";
		ram_buffer(9) := X"00A4182A";
		ram_buffer(10) := X"1460FFFD";
		ram_buffer(11) := X"24A50004";
		ram_buffer(12) := X"0C40007C";
		ram_buffer(13) := X"00000000";
		ram_buffer(14) := X"0840000E";
		ram_buffer(15) := X"23BDFF98";
		ram_buffer(16) := X"AFA10010";
		ram_buffer(17) := X"AFA20014";
		ram_buffer(18) := X"AFA30018";
		ram_buffer(19) := X"AFA4001C";
		ram_buffer(20) := X"AFA50020";
		ram_buffer(21) := X"AFA60024";
		ram_buffer(22) := X"AFA70028";
		ram_buffer(23) := X"AFA8002C";
		ram_buffer(24) := X"AFA90030";
		ram_buffer(25) := X"AFAA0034";
		ram_buffer(26) := X"AFAB0038";
		ram_buffer(27) := X"AFAC003C";
		ram_buffer(28) := X"AFAD0040";
		ram_buffer(29) := X"AFAE0044";
		ram_buffer(30) := X"AFAF0048";
		ram_buffer(31) := X"AFB8004C";
		ram_buffer(32) := X"AFB90050";
		ram_buffer(33) := X"AFBF0054";
		ram_buffer(34) := X"401A7000";
		ram_buffer(35) := X"235AFFFC";
		ram_buffer(36) := X"AFBA0058";
		ram_buffer(37) := X"0000D810";
		ram_buffer(38) := X"AFBB005C";
		ram_buffer(39) := X"0000D812";
		ram_buffer(40) := X"AFBB0060";
		ram_buffer(41) := X"0C4000C6";
		ram_buffer(42) := X"23A50000";
		ram_buffer(43) := X"8FA10010";
		ram_buffer(44) := X"8FA20014";
		ram_buffer(45) := X"8FA30018";
		ram_buffer(46) := X"8FA4001C";
		ram_buffer(47) := X"8FA50020";
		ram_buffer(48) := X"8FA60024";
		ram_buffer(49) := X"8FA70028";
		ram_buffer(50) := X"8FA8002C";
		ram_buffer(51) := X"8FA90030";
		ram_buffer(52) := X"8FAA0034";
		ram_buffer(53) := X"8FAB0038";
		ram_buffer(54) := X"8FAC003C";
		ram_buffer(55) := X"8FAD0040";
		ram_buffer(56) := X"8FAE0044";
		ram_buffer(57) := X"8FAF0048";
		ram_buffer(58) := X"8FB8004C";
		ram_buffer(59) := X"8FB90050";
		ram_buffer(60) := X"8FBF0054";
		ram_buffer(61) := X"8FBA0058";
		ram_buffer(62) := X"8FBB005C";
		ram_buffer(63) := X"03600011";
		ram_buffer(64) := X"8FBB0060";
		ram_buffer(65) := X"03600013";
		ram_buffer(66) := X"23BD0068";
		ram_buffer(67) := X"341B0001";
		ram_buffer(68) := X"03400008";
		ram_buffer(69) := X"409B6000";
		ram_buffer(70) := X"40026000";
		ram_buffer(71) := X"03E00008";
		ram_buffer(72) := X"40846000";
		ram_buffer(73) := X"3C050100";
		ram_buffer(74) := X"24A50150";
		ram_buffer(75) := X"8CA60000";
		ram_buffer(76) := X"AC06003C";
		ram_buffer(77) := X"8CA60004";
		ram_buffer(78) := X"AC060040";
		ram_buffer(79) := X"8CA60008";
		ram_buffer(80) := X"AC060044";
		ram_buffer(81) := X"8CA6000C";
		ram_buffer(82) := X"03E00008";
		ram_buffer(83) := X"AC060048";
		ram_buffer(84) := X"3C1A0100";
		ram_buffer(85) := X"375A003C";
		ram_buffer(86) := X"03400008";
		ram_buffer(87) := X"00000000";
		ram_buffer(88) := X"AC900000";
		ram_buffer(89) := X"AC910004";
		ram_buffer(90) := X"AC920008";
		ram_buffer(91) := X"AC93000C";
		ram_buffer(92) := X"AC940010";
		ram_buffer(93) := X"AC950014";
		ram_buffer(94) := X"AC960018";
		ram_buffer(95) := X"AC97001C";
		ram_buffer(96) := X"AC9E0020";
		ram_buffer(97) := X"AC9C0024";
		ram_buffer(98) := X"AC9D0028";
		ram_buffer(99) := X"AC9F002C";
		ram_buffer(100) := X"03E00008";
		ram_buffer(101) := X"34020000";
		ram_buffer(102) := X"8C900000";
		ram_buffer(103) := X"8C910004";
		ram_buffer(104) := X"8C920008";
		ram_buffer(105) := X"8C93000C";
		ram_buffer(106) := X"8C940010";
		ram_buffer(107) := X"8C950014";
		ram_buffer(108) := X"8C960018";
		ram_buffer(109) := X"8C97001C";
		ram_buffer(110) := X"8C9E0020";
		ram_buffer(111) := X"8C9C0024";
		ram_buffer(112) := X"8C9D0028";
		ram_buffer(113) := X"8C9F002C";
		ram_buffer(114) := X"03E00008";
		ram_buffer(115) := X"34A20000";
		ram_buffer(116) := X"00850019";
		ram_buffer(117) := X"00001012";
		ram_buffer(118) := X"00002010";
		ram_buffer(119) := X"03E00008";
		ram_buffer(120) := X"ACC40000";
		ram_buffer(121) := X"0000000C";
		ram_buffer(122) := X"03E00008";
		ram_buffer(123) := X"00000000";
		ram_buffer(124) := X"27BDFFE0";
		ram_buffer(125) := X"3C0244A0";
		ram_buffer(126) := X"AFB00014";
		ram_buffer(127) := X"3C100100";
		ram_buffer(128) := X"AE020A50";
		ram_buffer(129) := X"3C030100";
		ram_buffer(130) := X"3C020100";
		ram_buffer(131) := X"AFBF001C";
		ram_buffer(132) := X"AFB10018";
		ram_buffer(133) := X"24420A54";
		ram_buffer(134) := X"24630A94";
		ram_buffer(135) := X"24420008";
		ram_buffer(136) := X"1443FFFE";
		ram_buffer(137) := X"AC40FFF8";
		ram_buffer(138) := X"3C0244A2";
		ram_buffer(139) := X"AF828018";
		ram_buffer(140) := X"3C020100";
		ram_buffer(141) := X"26110A50";
		ram_buffer(142) := X"244202BC";
		ram_buffer(143) := X"3C050100";
		ram_buffer(144) := X"24A502E8";
		ram_buffer(145) := X"AE22000C";
		ram_buffer(146) := X"00002025";
		ram_buffer(147) := X"3C0244A4";
		ram_buffer(148) := X"AF82801C";
		ram_buffer(149) := X"0C4001E7";
		ram_buffer(150) := X"AE200010";
		ram_buffer(151) := X"3C020100";
		ram_buffer(152) := X"244202CC";
		ram_buffer(153) := X"AE22001C";
		ram_buffer(154) := X"0C400049";
		ram_buffer(155) := X"AE200020";
		ram_buffer(156) := X"0C400046";
		ram_buffer(157) := X"24040001";
		ram_buffer(158) := X"8E020A50";
		ram_buffer(159) := X"240300FF";
		ram_buffer(160) := X"AC430000";
		ram_buffer(161) := X"8F838018";
		ram_buffer(162) := X"24020001";
		ram_buffer(163) := X"AC620000";
		ram_buffer(164) := X"8F838018";
		ram_buffer(165) := X"3C040100";
		ram_buffer(166) := X"AC620008";
		ram_buffer(167) := X"0C4001EA";
		ram_buffer(168) := X"24840830";
		ram_buffer(169) := X"8FBF001C";
		ram_buffer(170) := X"8FB10018";
		ram_buffer(171) := X"8FB00014";
		ram_buffer(172) := X"00001025";
		ram_buffer(173) := X"03E00008";
		ram_buffer(174) := X"27BD0020";
		ram_buffer(175) := X"8F828018";
		ram_buffer(176) := X"24030003";
		ram_buffer(177) := X"03E00008";
		ram_buffer(178) := X"AC430000";
		ram_buffer(179) := X"8F82801C";
		ram_buffer(180) := X"00000000";
		ram_buffer(181) := X"8C430004";
		ram_buffer(182) := X"00000000";
		ram_buffer(183) := X"AC430008";
		ram_buffer(184) := X"03E00008";
		ram_buffer(185) := X"00000000";
		ram_buffer(186) := X"8F83801C";
		ram_buffer(187) := X"00000000";
		ram_buffer(188) := X"8C620000";
		ram_buffer(189) := X"00000000";
		ram_buffer(190) := X"30420002";
		ram_buffer(191) := X"10400003";
		ram_buffer(192) := X"00000000";
		ram_buffer(193) := X"03E00008";
		ram_buffer(194) := X"00000000";
		ram_buffer(195) := X"AC650008";
		ram_buffer(196) := X"1000FFF5";
		ram_buffer(197) := X"00000000";
		ram_buffer(198) := X"3C030100";
		ram_buffer(199) := X"8C620A50";
		ram_buffer(200) := X"27BDFFE0";
		ram_buffer(201) := X"8C420004";
		ram_buffer(202) := X"AFB10018";
		ram_buffer(203) := X"3C110100";
		ram_buffer(204) := X"AFB00014";
		ram_buffer(205) := X"AFBF001C";
		ram_buffer(206) := X"00608025";
		ram_buffer(207) := X"26310A54";
		ram_buffer(208) := X"2C430008";
		ram_buffer(209) := X"14600006";
		ram_buffer(210) := X"00000000";
		ram_buffer(211) := X"8FBF001C";
		ram_buffer(212) := X"8FB10018";
		ram_buffer(213) := X"8FB00014";
		ram_buffer(214) := X"03E00008";
		ram_buffer(215) := X"27BD0020";
		ram_buffer(216) := X"000210C0";
		ram_buffer(217) := X"02221021";
		ram_buffer(218) := X"8C430000";
		ram_buffer(219) := X"8C440004";
		ram_buffer(220) := X"0060F809";
		ram_buffer(221) := X"00000000";
		ram_buffer(222) := X"8E020A50";
		ram_buffer(223) := X"00000000";
		ram_buffer(224) := X"8C420004";
		ram_buffer(225) := X"1000FFEF";
		ram_buffer(226) := X"2C430008";
		ram_buffer(227) := X"10C0000D";
		ram_buffer(228) := X"00C53021";
		ram_buffer(229) := X"2402FFF0";
		ram_buffer(230) := X"00C21824";
		ram_buffer(231) := X"0066302B";
		ram_buffer(232) := X"00A22824";
		ram_buffer(233) := X"00063100";
		ram_buffer(234) := X"24620010";
		ram_buffer(235) := X"00463021";
		ram_buffer(236) := X"3C022000";
		ram_buffer(237) := X"00822021";
		ram_buffer(238) := X"2402FFF0";
		ram_buffer(239) := X"14C50003";
		ram_buffer(240) := X"00A21824";
		ram_buffer(241) := X"03E00008";
		ram_buffer(242) := X"00000000";
		ram_buffer(243) := X"AC830000";
		ram_buffer(244) := X"AC600000";
		ram_buffer(245) := X"1000FFF9";
		ram_buffer(246) := X"24A50010";
		ram_buffer(247) := X"24020001";
		ram_buffer(248) := X"14400002";
		ram_buffer(249) := X"0082001B";
		ram_buffer(250) := X"0007000D";
		ram_buffer(251) := X"00001812";
		ram_buffer(252) := X"0065182B";
		ram_buffer(253) := X"10600006";
		ram_buffer(254) := X"00450018";
		ram_buffer(255) := X"00004025";
		ram_buffer(256) := X"14400006";
		ram_buffer(257) := X"00000000";
		ram_buffer(258) := X"03E00008";
		ram_buffer(259) := X"A0E00000";
		ram_buffer(260) := X"00001012";
		ram_buffer(261) := X"1000FFF2";
		ram_buffer(262) := X"00000000";
		ram_buffer(263) := X"14400002";
		ram_buffer(264) := X"0082001B";
		ram_buffer(265) := X"0007000D";
		ram_buffer(266) := X"00002010";
		ram_buffer(267) := X"00004812";
		ram_buffer(268) := X"00000000";
		ram_buffer(269) := X"00000000";
		ram_buffer(270) := X"14A00002";
		ram_buffer(271) := X"0045001B";
		ram_buffer(272) := X"0007000D";
		ram_buffer(273) := X"00001012";
		ram_buffer(274) := X"15000005";
		ram_buffer(275) := X"292A000A";
		ram_buffer(276) := X"1D200004";
		ram_buffer(277) := X"24EB0001";
		ram_buffer(278) := X"1440FFE9";
		ram_buffer(279) := X"00000000";
		ram_buffer(280) := X"24EB0001";
		ram_buffer(281) := X"15400004";
		ram_buffer(282) := X"24030030";
		ram_buffer(283) := X"14C00002";
		ram_buffer(284) := X"24030037";
		ram_buffer(285) := X"24030057";
		ram_buffer(286) := X"00691821";
		ram_buffer(287) := X"A0E30000";
		ram_buffer(288) := X"25080001";
		ram_buffer(289) := X"1000FFDE";
		ram_buffer(290) := X"01603825";
		ram_buffer(291) := X"27BDFFD8";
		ram_buffer(292) := X"AFB40020";
		ram_buffer(293) := X"AFB3001C";
		ram_buffer(294) := X"AFB20018";
		ram_buffer(295) := X"AFB10014";
		ram_buffer(296) := X"AFBF0024";
		ram_buffer(297) := X"AFB00010";
		ram_buffer(298) := X"00809025";
		ram_buffer(299) := X"00A09825";
		ram_buffer(300) := X"8FB10038";
		ram_buffer(301) := X"10E00002";
		ram_buffer(302) := X"24140020";
		ram_buffer(303) := X"24140030";
		ram_buffer(304) := X"02201025";
		ram_buffer(305) := X"24420001";
		ram_buffer(306) := X"8043FFFF";
		ram_buffer(307) := X"00000000";
		ram_buffer(308) := X"14600009";
		ram_buffer(309) := X"00C08025";
		ram_buffer(310) := X"1A000009";
		ram_buffer(311) := X"02802825";
		ram_buffer(312) := X"0260F809";
		ram_buffer(313) := X"02402025";
		ram_buffer(314) := X"1000FFFB";
		ram_buffer(315) := X"2610FFFF";
		ram_buffer(316) := X"1000FFF4";
		ram_buffer(317) := X"24C6FFFF";
		ram_buffer(318) := X"1CC0FFFD";
		ram_buffer(319) := X"00000000";
		ram_buffer(320) := X"26310001";
		ram_buffer(321) := X"8225FFFF";
		ram_buffer(322) := X"00000000";
		ram_buffer(323) := X"14A00009";
		ram_buffer(324) := X"00000000";
		ram_buffer(325) := X"8FBF0024";
		ram_buffer(326) := X"8FB40020";
		ram_buffer(327) := X"8FB3001C";
		ram_buffer(328) := X"8FB20018";
		ram_buffer(329) := X"8FB10014";
		ram_buffer(330) := X"8FB00010";
		ram_buffer(331) := X"03E00008";
		ram_buffer(332) := X"27BD0028";
		ram_buffer(333) := X"0260F809";
		ram_buffer(334) := X"02402025";
		ram_buffer(335) := X"1000FFF1";
		ram_buffer(336) := X"26310001";
		ram_buffer(337) := X"8C820000";
		ram_buffer(338) := X"00000000";
		ram_buffer(339) := X"24430001";
		ram_buffer(340) := X"AC830000";
		ram_buffer(341) := X"03E00008";
		ram_buffer(342) := X"A0450000";
		ram_buffer(343) := X"27BDFFB8";
		ram_buffer(344) := X"AFB5003C";
		ram_buffer(345) := X"AFB40038";
		ram_buffer(346) := X"AFB30034";
		ram_buffer(347) := X"AFB20030";
		ram_buffer(348) := X"AFB1002C";
		ram_buffer(349) := X"AFB00028";
		ram_buffer(350) := X"AFBF0044";
		ram_buffer(351) := X"AFB60040";
		ram_buffer(352) := X"00809025";
		ram_buffer(353) := X"00A09825";
		ram_buffer(354) := X"00C08825";
		ram_buffer(355) := X"00E08025";
		ram_buffer(356) := X"24140025";
		ram_buffer(357) := X"24150030";
		ram_buffer(358) := X"82250000";
		ram_buffer(359) := X"00000000";
		ram_buffer(360) := X"10A00035";
		ram_buffer(361) := X"00000000";
		ram_buffer(362) := X"10B40006";
		ram_buffer(363) := X"00000000";
		ram_buffer(364) := X"26310001";
		ram_buffer(365) := X"0260F809";
		ram_buffer(366) := X"02402025";
		ram_buffer(367) := X"1000FFF6";
		ram_buffer(368) := X"00000000";
		ram_buffer(369) := X"82260001";
		ram_buffer(370) := X"00000000";
		ram_buffer(371) := X"10D50015";
		ram_buffer(372) := X"240D0001";
		ram_buffer(373) := X"26310002";
		ram_buffer(374) := X"00006825";
		ram_buffer(375) := X"24C2FFD0";
		ram_buffer(376) := X"304200FF";
		ram_buffer(377) := X"2C42000A";
		ram_buffer(378) := X"10400018";
		ram_buffer(379) := X"00006025";
		ram_buffer(380) := X"30C200FF";
		ram_buffer(381) := X"2443FFD0";
		ram_buffer(382) := X"2C63000A";
		ram_buffer(383) := X"1060000C";
		ram_buffer(384) := X"2443FF9F";
		ram_buffer(385) := X"24C3FFD0";
		ram_buffer(386) := X"000C1080";
		ram_buffer(387) := X"004C6021";
		ram_buffer(388) := X"000C6040";
		ram_buffer(389) := X"26310001";
		ram_buffer(390) := X"8226FFFF";
		ram_buffer(391) := X"1000FFF4";
		ram_buffer(392) := X"01836021";
		ram_buffer(393) := X"82260002";
		ram_buffer(394) := X"1000FFEC";
		ram_buffer(395) := X"26310003";
		ram_buffer(396) := X"2C630006";
		ram_buffer(397) := X"1060001A";
		ram_buffer(398) := X"2442FFBF";
		ram_buffer(399) := X"24C3FFA9";
		ram_buffer(400) := X"2862000B";
		ram_buffer(401) := X"1440FFF1";
		ram_buffer(402) := X"000C1080";
		ram_buffer(403) := X"24020063";
		ram_buffer(404) := X"10C20045";
		ram_buffer(405) := X"28C20064";
		ram_buffer(406) := X"10400016";
		ram_buffer(407) := X"24020073";
		ram_buffer(408) := X"10D4004C";
		ram_buffer(409) := X"24020058";
		ram_buffer(410) := X"10C20033";
		ram_buffer(411) := X"00000000";
		ram_buffer(412) := X"14C0FFC9";
		ram_buffer(413) := X"00000000";
		ram_buffer(414) := X"8FBF0044";
		ram_buffer(415) := X"8FB60040";
		ram_buffer(416) := X"8FB5003C";
		ram_buffer(417) := X"8FB40038";
		ram_buffer(418) := X"8FB30034";
		ram_buffer(419) := X"8FB20030";
		ram_buffer(420) := X"8FB1002C";
		ram_buffer(421) := X"8FB00028";
		ram_buffer(422) := X"03E00008";
		ram_buffer(423) := X"27BD0048";
		ram_buffer(424) := X"2C420006";
		ram_buffer(425) := X"1040FFEA";
		ram_buffer(426) := X"24020063";
		ram_buffer(427) := X"1000FFE4";
		ram_buffer(428) := X"24C3FFC9";
		ram_buffer(429) := X"10C20032";
		ram_buffer(430) := X"28C20074";
		ram_buffer(431) := X"10400019";
		ram_buffer(432) := X"24020075";
		ram_buffer(433) := X"24020064";
		ram_buffer(434) := X"14C2FFB3";
		ram_buffer(435) := X"26160004";
		ram_buffer(436) := X"8E040000";
		ram_buffer(437) := X"00000000";
		ram_buffer(438) := X"04810005";
		ram_buffer(439) := X"27A70018";
		ram_buffer(440) := X"2402002D";
		ram_buffer(441) := X"00042023";
		ram_buffer(442) := X"A3A20018";
		ram_buffer(443) := X"27A70019";
		ram_buffer(444) := X"00003025";
		ram_buffer(445) := X"2405000A";
		ram_buffer(446) := X"0C4000F7";
		ram_buffer(447) := X"00000000";
		ram_buffer(448) := X"27A20018";
		ram_buffer(449) := X"AFA20010";
		ram_buffer(450) := X"01A03825";
		ram_buffer(451) := X"01803025";
		ram_buffer(452) := X"02602825";
		ram_buffer(453) := X"0C400123";
		ram_buffer(454) := X"02402025";
		ram_buffer(455) := X"1000FF9E";
		ram_buffer(456) := X"02C08025";
		ram_buffer(457) := X"10C2000A";
		ram_buffer(458) := X"26160004";
		ram_buffer(459) := X"24020078";
		ram_buffer(460) := X"14C2FF99";
		ram_buffer(461) := X"00000000";
		ram_buffer(462) := X"38C60058";
		ram_buffer(463) := X"26160004";
		ram_buffer(464) := X"27A70018";
		ram_buffer(465) := X"2CC60001";
		ram_buffer(466) := X"10000004";
		ram_buffer(467) := X"24050010";
		ram_buffer(468) := X"27A70018";
		ram_buffer(469) := X"00003025";
		ram_buffer(470) := X"2405000A";
		ram_buffer(471) := X"8E040000";
		ram_buffer(472) := X"1000FFE5";
		ram_buffer(473) := X"00000000";
		ram_buffer(474) := X"82050003";
		ram_buffer(475) := X"02402025";
		ram_buffer(476) := X"0260F809";
		ram_buffer(477) := X"26160004";
		ram_buffer(478) := X"1000FF87";
		ram_buffer(479) := X"02C08025";
		ram_buffer(480) := X"8E020000";
		ram_buffer(481) := X"26160004";
		ram_buffer(482) := X"AFA20010";
		ram_buffer(483) := X"1000FFDF";
		ram_buffer(484) := X"00003825";
		ram_buffer(485) := X"1000FF87";
		ram_buffer(486) := X"24050025";
		ram_buffer(487) := X"AF858014";
		ram_buffer(488) := X"03E00008";
		ram_buffer(489) := X"AF848010";
		ram_buffer(490) := X"27BDFFE0";
		ram_buffer(491) := X"AFA50024";
		ram_buffer(492) := X"AFA60028";
		ram_buffer(493) := X"8F858014";
		ram_buffer(494) := X"00803025";
		ram_buffer(495) := X"8F848010";
		ram_buffer(496) := X"AFA7002C";
		ram_buffer(497) := X"27A70024";
		ram_buffer(498) := X"AFBF001C";
		ram_buffer(499) := X"0C400157";
		ram_buffer(500) := X"AFA70010";
		ram_buffer(501) := X"8FBF001C";
		ram_buffer(502) := X"00000000";
		ram_buffer(503) := X"03E00008";
		ram_buffer(504) := X"27BD0020";
		ram_buffer(505) := X"27BDFFE0";
		ram_buffer(506) := X"AFA60028";
		ram_buffer(507) := X"00A03025";
		ram_buffer(508) := X"3C050100";
		ram_buffer(509) := X"AFA40020";
		ram_buffer(510) := X"AFA7002C";
		ram_buffer(511) := X"27A40020";
		ram_buffer(512) := X"27A70028";
		ram_buffer(513) := X"24A50544";
		ram_buffer(514) := X"AFBF001C";
		ram_buffer(515) := X"0C400157";
		ram_buffer(516) := X"AFA70010";
		ram_buffer(517) := X"8FA20020";
		ram_buffer(518) := X"00000000";
		ram_buffer(519) := X"A0400000";
		ram_buffer(520) := X"8FBF001C";
		ram_buffer(521) := X"00000000";
		ram_buffer(522) := X"03E00008";
		ram_buffer(523) := X"27BD0020";
		ram_buffer(524) := X"48656C6C";
		ram_buffer(525) := X"6F20576F";
		ram_buffer(526) := X"726C6421";
		ram_buffer(527) := X"0A0D0000";
		ram_buffer(528) := X"00000000";
		ram_buffer(529) := X"00000000";
		ram_buffer(530) := X"00000000";
		ram_buffer(531) := X"00000000";
		ram_buffer(532) := X"00000000";
		ram_buffer(533) := X"00000000";
		ram_buffer(534) := X"00000000";
		ram_buffer(535) := X"00000000";
		ram_buffer(536) := X"00000000";
		ram_buffer(537) := X"00000000";
		ram_buffer(538) := X"00000000";
		ram_buffer(539) := X"00000000";
		ram_buffer(540) := X"00000000";
		ram_buffer(541) := X"00000000";
		ram_buffer(542) := X"00000000";
		ram_buffer(543) := X"00000000";
		ram_buffer(544) := X"00000000";
		ram_buffer(545) := X"00000000";
		ram_buffer(546) := X"00000000";
		ram_buffer(547) := X"00000000";
		ram_buffer(548) := X"00000000";
		ram_buffer(549) := X"00000000";
		ram_buffer(550) := X"00000000";
		ram_buffer(551) := X"00000000";
		ram_buffer(552) := X"00000000";
		ram_buffer(553) := X"00000000";
		ram_buffer(554) := X"00000000";
		ram_buffer(555) := X"00000000";
		ram_buffer(556) := X"00000000";
		ram_buffer(557) := X"00000000";
		ram_buffer(558) := X"00000000";
		ram_buffer(559) := X"00000000";
		ram_buffer(560) := X"00000000";
		ram_buffer(561) := X"00000000";
		ram_buffer(562) := X"00000000";
		ram_buffer(563) := X"00000000";
		ram_buffer(564) := X"00000000";
		ram_buffer(565) := X"00000000";
		ram_buffer(566) := X"00000000";
		ram_buffer(567) := X"00000000";
		ram_buffer(568) := X"00000000";
		ram_buffer(569) := X"00000000";
		ram_buffer(570) := X"00000000";
		ram_buffer(571) := X"00000000";
		ram_buffer(572) := X"00000000";
		ram_buffer(573) := X"00000000";
		ram_buffer(574) := X"00000000";
		ram_buffer(575) := X"00000000";
		ram_buffer(576) := X"00000000";
		ram_buffer(577) := X"00000000";
		ram_buffer(578) := X"00000000";
		ram_buffer(579) := X"00000000";
		ram_buffer(580) := X"00000000";
		ram_buffer(581) := X"00000000";
		ram_buffer(582) := X"00000000";
		ram_buffer(583) := X"00000000";
		ram_buffer(584) := X"00000000";
		ram_buffer(585) := X"00000000";
		ram_buffer(586) := X"00000000";
		ram_buffer(587) := X"00000000";
		ram_buffer(588) := X"00000000";
		ram_buffer(589) := X"00000000";
		ram_buffer(590) := X"00000000";
		ram_buffer(591) := X"00000000";
		ram_buffer(592) := X"00000000";
		ram_buffer(593) := X"00000000";
		ram_buffer(594) := X"00000000";
		ram_buffer(595) := X"00000000";
		ram_buffer(596) := X"00000000";
		ram_buffer(597) := X"00000000";
		ram_buffer(598) := X"00000000";
		ram_buffer(599) := X"00000000";
		ram_buffer(600) := X"00000000";
		ram_buffer(601) := X"00000000";
		ram_buffer(602) := X"00000000";
		ram_buffer(603) := X"00000000";
		ram_buffer(604) := X"00000000";
		ram_buffer(605) := X"00000000";
		ram_buffer(606) := X"00000000";
		ram_buffer(607) := X"00000000";
		ram_buffer(608) := X"00000000";
		ram_buffer(609) := X"00000000";
		ram_buffer(610) := X"00000000";
		ram_buffer(611) := X"00000000";
		ram_buffer(612) := X"00000000";
		ram_buffer(613) := X"00000000";
		ram_buffer(614) := X"00000000";
		ram_buffer(615) := X"00000000";
		ram_buffer(616) := X"00000000";
		ram_buffer(617) := X"00000000";
		ram_buffer(618) := X"00000000";
		ram_buffer(619) := X"00000000";
		ram_buffer(620) := X"00000000";
		ram_buffer(621) := X"00000000";
		ram_buffer(622) := X"00000000";
		ram_buffer(623) := X"00000000";
		ram_buffer(624) := X"00000000";
		ram_buffer(625) := X"00000000";
		ram_buffer(626) := X"00000000";
		ram_buffer(627) := X"00000000";
		ram_buffer(628) := X"00000000";
		ram_buffer(629) := X"00000000";
		ram_buffer(630) := X"00000000";
		ram_buffer(631) := X"00000000";
		ram_buffer(632) := X"00000000";
		ram_buffer(633) := X"00000000";
		ram_buffer(634) := X"00000000";
		ram_buffer(635) := X"00000000";
		ram_buffer(636) := X"00000000";
		ram_buffer(637) := X"00000000";
		ram_buffer(638) := X"00000000";
		ram_buffer(639) := X"00000000";
		ram_buffer(640) := X"00000000";
		ram_buffer(641) := X"00000000";
		ram_buffer(642) := X"00000000";
		ram_buffer(643) := X"00000000";
		ram_buffer(644) := X"00000000";
		ram_buffer(645) := X"00000000";
		ram_buffer(646) := X"00000000";
		ram_buffer(647) := X"00000000";
		ram_buffer(648) := X"00000000";
		ram_buffer(649) := X"00000000";
		ram_buffer(650) := X"00000000";
		ram_buffer(651) := X"00000000";
		ram_buffer(652) := X"00000000";
		ram_buffer(653) := X"00000000";
		ram_buffer(654) := X"00000000";
		ram_buffer(655) := X"00000000";
		ram_buffer(656) := X"00000000";
		ram_buffer(657) := X"00000000";
		ram_buffer(658) := X"00000000";
		ram_buffer(659) := X"00000000";
		ram_buffer(660) := X"00000000";
		ram_buffer(661) := X"00000000";
		ram_buffer(662) := X"00000000";
		ram_buffer(663) := X"00000000";
		ram_buffer(664) := X"00000000";
		ram_buffer(665) := X"00000000";
		ram_buffer(666) := X"00000000";
		ram_buffer(667) := X"00000000";
		ram_buffer(668) := X"00000000";
		ram_buffer(669) := X"00000000";
		ram_buffer(670) := X"00000000";
		ram_buffer(671) := X"00000000";
		ram_buffer(672) := X"00000000";
		ram_buffer(673) := X"00000000";
		ram_buffer(674) := X"00000000";
		ram_buffer(675) := X"00000000";
		ram_buffer(676) := X"00000000";
		ram_buffer(677) := X"00000000";
		ram_buffer(678) := X"00000000";
		ram_buffer(679) := X"00000000";
		ram_buffer(680) := X"00000000";
		ram_buffer(681) := X"00000000";
		ram_buffer(682) := X"00000000";
		ram_buffer(683) := X"00000000";
		ram_buffer(684) := X"00000000";
		ram_buffer(685) := X"00000000";
		ram_buffer(686) := X"00000000";
		ram_buffer(687) := X"00000000";
		ram_buffer(688) := X"00000000";
		ram_buffer(689) := X"00000000";
		ram_buffer(690) := X"00000000";
		ram_buffer(691) := X"00000000";
		ram_buffer(692) := X"00000000";
		ram_buffer(693) := X"00000000";
		ram_buffer(694) := X"00000000";
		ram_buffer(695) := X"00000000";
		ram_buffer(696) := X"00000000";
		ram_buffer(697) := X"00000000";
		ram_buffer(698) := X"00000000";
		ram_buffer(699) := X"00000000";
		ram_buffer(700) := X"00000000";
		ram_buffer(701) := X"00000000";
		ram_buffer(702) := X"00000000";
		ram_buffer(703) := X"00000000";
		ram_buffer(704) := X"00000100";
		ram_buffer(705) := X"01010001";
		ram_buffer(706) := X"00000000";
		ram_buffer(707) := X"00000000";
		ram_buffer(708) := X"00000000";
		ram_buffer(709) := X"00000000";
		return ram_buffer;
	end;
end;
