library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.numeric_std.all;

package plasoc_gpio_pack is

end;

package body plasoc_gpio_pack is

end;